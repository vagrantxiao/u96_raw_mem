`timescale 1 ns / 1 ps

(* CORE_GENERATION_INFO = "vadd_bw_vadd_bw,hls_ip_2022_2,{HLS_INPUT_TYPE=cxx,HLS_INPUT_FLOAT=0,HLS_INPUT_FIXED=0,HLS_INPUT_PART=xcu50-fsvh2104-2-e,HLS_INPUT_CLOCK=3.330000,HLS_INPUT_ARCH=others,HLS_SYN_CLOCK=1.000000,HLS_SYN_LAT=0,HLS_SYN_TPT=none,HLS_SYN_MEM=0,HLS_SYN_DSP=0,HLS_SYN_FF=2066,HLS_SYN_LUT=3752,HLS_VERSION=2022_2}" *)


module vadd_bw
(
  s_axi_control_AWVALID,
  s_axi_control_AWREADY,
  s_axi_control_AWADDR,
  s_axi_control_WVALID,
  s_axi_control_WREADY,
  s_axi_control_WDATA,
  s_axi_control_WSTRB,
  s_axi_control_ARVALID,
  s_axi_control_ARREADY,
  s_axi_control_ARADDR,
  s_axi_control_RVALID,
  s_axi_control_RREADY,
  s_axi_control_RDATA,
  s_axi_control_RRESP,
  s_axi_control_BVALID,
  s_axi_control_BREADY,
  s_axi_control_BRESP,
  ap_clk,
  ap_rst_n,
  interrupt,
  m_axi_rmem0_ARADDR,
  m_axi_rmem0_ARBURST,
  m_axi_rmem0_ARCACHE,
  m_axi_rmem0_ARID,
  m_axi_rmem0_ARLEN,
  m_axi_rmem0_ARLOCK,
  m_axi_rmem0_ARPROT,
  m_axi_rmem0_ARQOS,
  m_axi_rmem0_ARREADY,
  m_axi_rmem0_ARSIZE,
  m_axi_rmem0_ARVALID,
  m_axi_rmem0_AWADDR,
  m_axi_rmem0_AWBURST,
  m_axi_rmem0_AWCACHE,
  m_axi_rmem0_AWID,
  m_axi_rmem0_AWLEN,
  m_axi_rmem0_AWLOCK,
  m_axi_rmem0_AWPROT,
  m_axi_rmem0_AWQOS,
  m_axi_rmem0_AWREADY,
  m_axi_rmem0_AWSIZE,
  m_axi_rmem0_AWVALID,
  m_axi_rmem0_BID,
  m_axi_rmem0_BREADY,
  m_axi_rmem0_BRESP,
  m_axi_rmem0_BVALID,
  m_axi_rmem0_RDATA,
  m_axi_rmem0_RID,
  m_axi_rmem0_RLAST,
  m_axi_rmem0_RREADY,
  m_axi_rmem0_RRESP,
  m_axi_rmem0_RVALID,
  m_axi_rmem0_WDATA,
  m_axi_rmem0_WLAST,
  m_axi_rmem0_WREADY,
  m_axi_rmem0_WSTRB,
  m_axi_rmem0_WVALID,
  m_axi_rmem1_ARADDR,
  m_axi_rmem1_ARBURST,
  m_axi_rmem1_ARCACHE,
  m_axi_rmem1_ARID,
  m_axi_rmem1_ARLEN,
  m_axi_rmem1_ARLOCK,
  m_axi_rmem1_ARPROT,
  m_axi_rmem1_ARQOS,
  m_axi_rmem1_ARREADY,
  m_axi_rmem1_ARSIZE,
  m_axi_rmem1_ARVALID,
  m_axi_rmem1_AWADDR,
  m_axi_rmem1_AWBURST,
  m_axi_rmem1_AWCACHE,
  m_axi_rmem1_AWID,
  m_axi_rmem1_AWLEN,
  m_axi_rmem1_AWLOCK,
  m_axi_rmem1_AWPROT,
  m_axi_rmem1_AWQOS,
  m_axi_rmem1_AWREADY,
  m_axi_rmem1_AWSIZE,
  m_axi_rmem1_AWVALID,
  m_axi_rmem1_BID,
  m_axi_rmem1_BREADY,
  m_axi_rmem1_BRESP,
  m_axi_rmem1_BVALID,
  m_axi_rmem1_RDATA,
  m_axi_rmem1_RID,
  m_axi_rmem1_RLAST,
  m_axi_rmem1_RREADY,
  m_axi_rmem1_RRESP,
  m_axi_rmem1_RVALID,
  m_axi_rmem1_WDATA,
  m_axi_rmem1_WLAST,
  m_axi_rmem1_WREADY,
  m_axi_rmem1_WSTRB,
  m_axi_rmem1_WVALID,
  m_axi_rmem2_ARADDR,
  m_axi_rmem2_ARBURST,
  m_axi_rmem2_ARCACHE,
  m_axi_rmem2_ARID,
  m_axi_rmem2_ARLEN,
  m_axi_rmem2_ARLOCK,
  m_axi_rmem2_ARPROT,
  m_axi_rmem2_ARQOS,
  m_axi_rmem2_ARREADY,
  m_axi_rmem2_ARSIZE,
  m_axi_rmem2_ARVALID,
  m_axi_rmem2_AWADDR,
  m_axi_rmem2_AWBURST,
  m_axi_rmem2_AWCACHE,
  m_axi_rmem2_AWID,
  m_axi_rmem2_AWLEN,
  m_axi_rmem2_AWLOCK,
  m_axi_rmem2_AWPROT,
  m_axi_rmem2_AWQOS,
  m_axi_rmem2_AWREADY,
  m_axi_rmem2_AWSIZE,
  m_axi_rmem2_AWVALID,
  m_axi_rmem2_BID,
  m_axi_rmem2_BREADY,
  m_axi_rmem2_BRESP,
  m_axi_rmem2_BVALID,
  m_axi_rmem2_RDATA,
  m_axi_rmem2_RID,
  m_axi_rmem2_RLAST,
  m_axi_rmem2_RREADY,
  m_axi_rmem2_RRESP,
  m_axi_rmem2_RVALID,
  m_axi_rmem2_WDATA,
  m_axi_rmem2_WLAST,
  m_axi_rmem2_WREADY,
  m_axi_rmem2_WSTRB,
  m_axi_rmem2_WVALID,
  m_axi_rmem3_ARADDR,
  m_axi_rmem3_ARBURST,
  m_axi_rmem3_ARCACHE,
  m_axi_rmem3_ARID,
  m_axi_rmem3_ARLEN,
  m_axi_rmem3_ARLOCK,
  m_axi_rmem3_ARPROT,
  m_axi_rmem3_ARQOS,
  m_axi_rmem3_ARREADY,
  m_axi_rmem3_ARSIZE,
  m_axi_rmem3_ARVALID,
  m_axi_rmem3_AWADDR,
  m_axi_rmem3_AWBURST,
  m_axi_rmem3_AWCACHE,
  m_axi_rmem3_AWID,
  m_axi_rmem3_AWLEN,
  m_axi_rmem3_AWLOCK,
  m_axi_rmem3_AWPROT,
  m_axi_rmem3_AWQOS,
  m_axi_rmem3_AWREADY,
  m_axi_rmem3_AWSIZE,
  m_axi_rmem3_AWVALID,
  m_axi_rmem3_BID,
  m_axi_rmem3_BREADY,
  m_axi_rmem3_BRESP,
  m_axi_rmem3_BVALID,
  m_axi_rmem3_RDATA,
  m_axi_rmem3_RID,
  m_axi_rmem3_RLAST,
  m_axi_rmem3_RREADY,
  m_axi_rmem3_RRESP,
  m_axi_rmem3_RVALID,
  m_axi_rmem3_WDATA,
  m_axi_rmem3_WLAST,
  m_axi_rmem3_WREADY,
  m_axi_rmem3_WSTRB,
  m_axi_rmem3_WVALID,
  m_axi_rmem4_ARADDR,
  m_axi_rmem4_ARBURST,
  m_axi_rmem4_ARCACHE,
  m_axi_rmem4_ARID,
  m_axi_rmem4_ARLEN,
  m_axi_rmem4_ARLOCK,
  m_axi_rmem4_ARPROT,
  m_axi_rmem4_ARQOS,
  m_axi_rmem4_ARREADY,
  m_axi_rmem4_ARSIZE,
  m_axi_rmem4_ARVALID,
  m_axi_rmem4_AWADDR,
  m_axi_rmem4_AWBURST,
  m_axi_rmem4_AWCACHE,
  m_axi_rmem4_AWID,
  m_axi_rmem4_AWLEN,
  m_axi_rmem4_AWLOCK,
  m_axi_rmem4_AWPROT,
  m_axi_rmem4_AWQOS,
  m_axi_rmem4_AWREADY,
  m_axi_rmem4_AWSIZE,
  m_axi_rmem4_AWVALID,
  m_axi_rmem4_BID,
  m_axi_rmem4_BREADY,
  m_axi_rmem4_BRESP,
  m_axi_rmem4_BVALID,
  m_axi_rmem4_RDATA,
  m_axi_rmem4_RID,
  m_axi_rmem4_RLAST,
  m_axi_rmem4_RREADY,
  m_axi_rmem4_RRESP,
  m_axi_rmem4_RVALID,
  m_axi_rmem4_WDATA,
  m_axi_rmem4_WLAST,
  m_axi_rmem4_WREADY,
  m_axi_rmem4_WSTRB,
  m_axi_rmem4_WVALID,
  m_axi_rmem5_ARADDR,
  m_axi_rmem5_ARBURST,
  m_axi_rmem5_ARCACHE,
  m_axi_rmem5_ARID,
  m_axi_rmem5_ARLEN,
  m_axi_rmem5_ARLOCK,
  m_axi_rmem5_ARPROT,
  m_axi_rmem5_ARQOS,
  m_axi_rmem5_ARREADY,
  m_axi_rmem5_ARSIZE,
  m_axi_rmem5_ARVALID,
  m_axi_rmem5_AWADDR,
  m_axi_rmem5_AWBURST,
  m_axi_rmem5_AWCACHE,
  m_axi_rmem5_AWID,
  m_axi_rmem5_AWLEN,
  m_axi_rmem5_AWLOCK,
  m_axi_rmem5_AWPROT,
  m_axi_rmem5_AWQOS,
  m_axi_rmem5_AWREADY,
  m_axi_rmem5_AWSIZE,
  m_axi_rmem5_AWVALID,
  m_axi_rmem5_BID,
  m_axi_rmem5_BREADY,
  m_axi_rmem5_BRESP,
  m_axi_rmem5_BVALID,
  m_axi_rmem5_RDATA,
  m_axi_rmem5_RID,
  m_axi_rmem5_RLAST,
  m_axi_rmem5_RREADY,
  m_axi_rmem5_RRESP,
  m_axi_rmem5_RVALID,
  m_axi_rmem5_WDATA,
  m_axi_rmem5_WLAST,
  m_axi_rmem5_WREADY,
  m_axi_rmem5_WSTRB,
  m_axi_rmem5_WVALID,
  m_axi_rmem6_ARADDR,
  m_axi_rmem6_ARBURST,
  m_axi_rmem6_ARCACHE,
  m_axi_rmem6_ARID,
  m_axi_rmem6_ARLEN,
  m_axi_rmem6_ARLOCK,
  m_axi_rmem6_ARPROT,
  m_axi_rmem6_ARQOS,
  m_axi_rmem6_ARREADY,
  m_axi_rmem6_ARSIZE,
  m_axi_rmem6_ARVALID,
  m_axi_rmem6_AWADDR,
  m_axi_rmem6_AWBURST,
  m_axi_rmem6_AWCACHE,
  m_axi_rmem6_AWID,
  m_axi_rmem6_AWLEN,
  m_axi_rmem6_AWLOCK,
  m_axi_rmem6_AWPROT,
  m_axi_rmem6_AWQOS,
  m_axi_rmem6_AWREADY,
  m_axi_rmem6_AWSIZE,
  m_axi_rmem6_AWVALID,
  m_axi_rmem6_BID,
  m_axi_rmem6_BREADY,
  m_axi_rmem6_BRESP,
  m_axi_rmem6_BVALID,
  m_axi_rmem6_RDATA,
  m_axi_rmem6_RID,
  m_axi_rmem6_RLAST,
  m_axi_rmem6_RREADY,
  m_axi_rmem6_RRESP,
  m_axi_rmem6_RVALID,
  m_axi_rmem6_WDATA,
  m_axi_rmem6_WLAST,
  m_axi_rmem6_WREADY,
  m_axi_rmem6_WSTRB,
  m_axi_rmem6_WVALID,
  m_axi_rmem7_ARADDR,
  m_axi_rmem7_ARBURST,
  m_axi_rmem7_ARCACHE,
  m_axi_rmem7_ARID,
  m_axi_rmem7_ARLEN,
  m_axi_rmem7_ARLOCK,
  m_axi_rmem7_ARPROT,
  m_axi_rmem7_ARQOS,
  m_axi_rmem7_ARREADY,
  m_axi_rmem7_ARSIZE,
  m_axi_rmem7_ARVALID,
  m_axi_rmem7_AWADDR,
  m_axi_rmem7_AWBURST,
  m_axi_rmem7_AWCACHE,
  m_axi_rmem7_AWID,
  m_axi_rmem7_AWLEN,
  m_axi_rmem7_AWLOCK,
  m_axi_rmem7_AWPROT,
  m_axi_rmem7_AWQOS,
  m_axi_rmem7_AWREADY,
  m_axi_rmem7_AWSIZE,
  m_axi_rmem7_AWVALID,
  m_axi_rmem7_BID,
  m_axi_rmem7_BREADY,
  m_axi_rmem7_BRESP,
  m_axi_rmem7_BVALID,
  m_axi_rmem7_RDATA,
  m_axi_rmem7_RID,
  m_axi_rmem7_RLAST,
  m_axi_rmem7_RREADY,
  m_axi_rmem7_RRESP,
  m_axi_rmem7_RVALID,
  m_axi_rmem7_WDATA,
  m_axi_rmem7_WLAST,
  m_axi_rmem7_WREADY,
  m_axi_rmem7_WSTRB,
  m_axi_rmem7_WVALID,
  m_axi_rmem8_ARADDR,
  m_axi_rmem8_ARBURST,
  m_axi_rmem8_ARCACHE,
  m_axi_rmem8_ARID,
  m_axi_rmem8_ARLEN,
  m_axi_rmem8_ARLOCK,
  m_axi_rmem8_ARPROT,
  m_axi_rmem8_ARQOS,
  m_axi_rmem8_ARREADY,
  m_axi_rmem8_ARSIZE,
  m_axi_rmem8_ARVALID,
  m_axi_rmem8_AWADDR,
  m_axi_rmem8_AWBURST,
  m_axi_rmem8_AWCACHE,
  m_axi_rmem8_AWID,
  m_axi_rmem8_AWLEN,
  m_axi_rmem8_AWLOCK,
  m_axi_rmem8_AWPROT,
  m_axi_rmem8_AWQOS,
  m_axi_rmem8_AWREADY,
  m_axi_rmem8_AWSIZE,
  m_axi_rmem8_AWVALID,
  m_axi_rmem8_BID,
  m_axi_rmem8_BREADY,
  m_axi_rmem8_BRESP,
  m_axi_rmem8_BVALID,
  m_axi_rmem8_RDATA,
  m_axi_rmem8_RID,
  m_axi_rmem8_RLAST,
  m_axi_rmem8_RREADY,
  m_axi_rmem8_RRESP,
  m_axi_rmem8_RVALID,
  m_axi_rmem8_WDATA,
  m_axi_rmem8_WLAST,
  m_axi_rmem8_WREADY,
  m_axi_rmem8_WSTRB,
  m_axi_rmem8_WVALID,
  m_axi_rmem9_ARADDR,
  m_axi_rmem9_ARBURST,
  m_axi_rmem9_ARCACHE,
  m_axi_rmem9_ARID,
  m_axi_rmem9_ARLEN,
  m_axi_rmem9_ARLOCK,
  m_axi_rmem9_ARPROT,
  m_axi_rmem9_ARQOS,
  m_axi_rmem9_ARREADY,
  m_axi_rmem9_ARSIZE,
  m_axi_rmem9_ARVALID,
  m_axi_rmem9_AWADDR,
  m_axi_rmem9_AWBURST,
  m_axi_rmem9_AWCACHE,
  m_axi_rmem9_AWID,
  m_axi_rmem9_AWLEN,
  m_axi_rmem9_AWLOCK,
  m_axi_rmem9_AWPROT,
  m_axi_rmem9_AWQOS,
  m_axi_rmem9_AWREADY,
  m_axi_rmem9_AWSIZE,
  m_axi_rmem9_AWVALID,
  m_axi_rmem9_BID,
  m_axi_rmem9_BREADY,
  m_axi_rmem9_BRESP,
  m_axi_rmem9_BVALID,
  m_axi_rmem9_RDATA,
  m_axi_rmem9_RID,
  m_axi_rmem9_RLAST,
  m_axi_rmem9_RREADY,
  m_axi_rmem9_RRESP,
  m_axi_rmem9_RVALID,
  m_axi_rmem9_WDATA,
  m_axi_rmem9_WLAST,
  m_axi_rmem9_WREADY,
  m_axi_rmem9_WSTRB,
  m_axi_rmem9_WVALID,
  m_axi_rmem10_ARADDR,
  m_axi_rmem10_ARBURST,
  m_axi_rmem10_ARCACHE,
  m_axi_rmem10_ARID,
  m_axi_rmem10_ARLEN,
  m_axi_rmem10_ARLOCK,
  m_axi_rmem10_ARPROT,
  m_axi_rmem10_ARQOS,
  m_axi_rmem10_ARREADY,
  m_axi_rmem10_ARSIZE,
  m_axi_rmem10_ARVALID,
  m_axi_rmem10_AWADDR,
  m_axi_rmem10_AWBURST,
  m_axi_rmem10_AWCACHE,
  m_axi_rmem10_AWID,
  m_axi_rmem10_AWLEN,
  m_axi_rmem10_AWLOCK,
  m_axi_rmem10_AWPROT,
  m_axi_rmem10_AWQOS,
  m_axi_rmem10_AWREADY,
  m_axi_rmem10_AWSIZE,
  m_axi_rmem10_AWVALID,
  m_axi_rmem10_BID,
  m_axi_rmem10_BREADY,
  m_axi_rmem10_BRESP,
  m_axi_rmem10_BVALID,
  m_axi_rmem10_RDATA,
  m_axi_rmem10_RID,
  m_axi_rmem10_RLAST,
  m_axi_rmem10_RREADY,
  m_axi_rmem10_RRESP,
  m_axi_rmem10_RVALID,
  m_axi_rmem10_WDATA,
  m_axi_rmem10_WLAST,
  m_axi_rmem10_WREADY,
  m_axi_rmem10_WSTRB,
  m_axi_rmem10_WVALID,
  m_axi_rmem11_ARADDR,
  m_axi_rmem11_ARBURST,
  m_axi_rmem11_ARCACHE,
  m_axi_rmem11_ARID,
  m_axi_rmem11_ARLEN,
  m_axi_rmem11_ARLOCK,
  m_axi_rmem11_ARPROT,
  m_axi_rmem11_ARQOS,
  m_axi_rmem11_ARREADY,
  m_axi_rmem11_ARSIZE,
  m_axi_rmem11_ARVALID,
  m_axi_rmem11_AWADDR,
  m_axi_rmem11_AWBURST,
  m_axi_rmem11_AWCACHE,
  m_axi_rmem11_AWID,
  m_axi_rmem11_AWLEN,
  m_axi_rmem11_AWLOCK,
  m_axi_rmem11_AWPROT,
  m_axi_rmem11_AWQOS,
  m_axi_rmem11_AWREADY,
  m_axi_rmem11_AWSIZE,
  m_axi_rmem11_AWVALID,
  m_axi_rmem11_BID,
  m_axi_rmem11_BREADY,
  m_axi_rmem11_BRESP,
  m_axi_rmem11_BVALID,
  m_axi_rmem11_RDATA,
  m_axi_rmem11_RID,
  m_axi_rmem11_RLAST,
  m_axi_rmem11_RREADY,
  m_axi_rmem11_RRESP,
  m_axi_rmem11_RVALID,
  m_axi_rmem11_WDATA,
  m_axi_rmem11_WLAST,
  m_axi_rmem11_WREADY,
  m_axi_rmem11_WSTRB,
  m_axi_rmem11_WVALID,
  m_axi_rmem12_ARADDR,
  m_axi_rmem12_ARBURST,
  m_axi_rmem12_ARCACHE,
  m_axi_rmem12_ARID,
  m_axi_rmem12_ARLEN,
  m_axi_rmem12_ARLOCK,
  m_axi_rmem12_ARPROT,
  m_axi_rmem12_ARQOS,
  m_axi_rmem12_ARREADY,
  m_axi_rmem12_ARSIZE,
  m_axi_rmem12_ARVALID,
  m_axi_rmem12_AWADDR,
  m_axi_rmem12_AWBURST,
  m_axi_rmem12_AWCACHE,
  m_axi_rmem12_AWID,
  m_axi_rmem12_AWLEN,
  m_axi_rmem12_AWLOCK,
  m_axi_rmem12_AWPROT,
  m_axi_rmem12_AWQOS,
  m_axi_rmem12_AWREADY,
  m_axi_rmem12_AWSIZE,
  m_axi_rmem12_AWVALID,
  m_axi_rmem12_BID,
  m_axi_rmem12_BREADY,
  m_axi_rmem12_BRESP,
  m_axi_rmem12_BVALID,
  m_axi_rmem12_RDATA,
  m_axi_rmem12_RID,
  m_axi_rmem12_RLAST,
  m_axi_rmem12_RREADY,
  m_axi_rmem12_RRESP,
  m_axi_rmem12_RVALID,
  m_axi_rmem12_WDATA,
  m_axi_rmem12_WLAST,
  m_axi_rmem12_WREADY,
  m_axi_rmem12_WSTRB,
  m_axi_rmem12_WVALID,
  m_axi_rmem13_ARADDR,
  m_axi_rmem13_ARBURST,
  m_axi_rmem13_ARCACHE,
  m_axi_rmem13_ARID,
  m_axi_rmem13_ARLEN,
  m_axi_rmem13_ARLOCK,
  m_axi_rmem13_ARPROT,
  m_axi_rmem13_ARQOS,
  m_axi_rmem13_ARREADY,
  m_axi_rmem13_ARSIZE,
  m_axi_rmem13_ARVALID,
  m_axi_rmem13_AWADDR,
  m_axi_rmem13_AWBURST,
  m_axi_rmem13_AWCACHE,
  m_axi_rmem13_AWID,
  m_axi_rmem13_AWLEN,
  m_axi_rmem13_AWLOCK,
  m_axi_rmem13_AWPROT,
  m_axi_rmem13_AWQOS,
  m_axi_rmem13_AWREADY,
  m_axi_rmem13_AWSIZE,
  m_axi_rmem13_AWVALID,
  m_axi_rmem13_BID,
  m_axi_rmem13_BREADY,
  m_axi_rmem13_BRESP,
  m_axi_rmem13_BVALID,
  m_axi_rmem13_RDATA,
  m_axi_rmem13_RID,
  m_axi_rmem13_RLAST,
  m_axi_rmem13_RREADY,
  m_axi_rmem13_RRESP,
  m_axi_rmem13_RVALID,
  m_axi_rmem13_WDATA,
  m_axi_rmem13_WLAST,
  m_axi_rmem13_WREADY,
  m_axi_rmem13_WSTRB,
  m_axi_rmem13_WVALID,
  m_axi_rmem14_ARADDR,
  m_axi_rmem14_ARBURST,
  m_axi_rmem14_ARCACHE,
  m_axi_rmem14_ARID,
  m_axi_rmem14_ARLEN,
  m_axi_rmem14_ARLOCK,
  m_axi_rmem14_ARPROT,
  m_axi_rmem14_ARQOS,
  m_axi_rmem14_ARREADY,
  m_axi_rmem14_ARSIZE,
  m_axi_rmem14_ARVALID,
  m_axi_rmem14_AWADDR,
  m_axi_rmem14_AWBURST,
  m_axi_rmem14_AWCACHE,
  m_axi_rmem14_AWID,
  m_axi_rmem14_AWLEN,
  m_axi_rmem14_AWLOCK,
  m_axi_rmem14_AWPROT,
  m_axi_rmem14_AWQOS,
  m_axi_rmem14_AWREADY,
  m_axi_rmem14_AWSIZE,
  m_axi_rmem14_AWVALID,
  m_axi_rmem14_BID,
  m_axi_rmem14_BREADY,
  m_axi_rmem14_BRESP,
  m_axi_rmem14_BVALID,
  m_axi_rmem14_RDATA,
  m_axi_rmem14_RID,
  m_axi_rmem14_RLAST,
  m_axi_rmem14_RREADY,
  m_axi_rmem14_RRESP,
  m_axi_rmem14_RVALID,
  m_axi_rmem14_WDATA,
  m_axi_rmem14_WLAST,
  m_axi_rmem14_WREADY,
  m_axi_rmem14_WSTRB,
  m_axi_rmem14_WVALID,
  m_axi_rmem15_ARADDR,
  m_axi_rmem15_ARBURST,
  m_axi_rmem15_ARCACHE,
  m_axi_rmem15_ARID,
  m_axi_rmem15_ARLEN,
  m_axi_rmem15_ARLOCK,
  m_axi_rmem15_ARPROT,
  m_axi_rmem15_ARQOS,
  m_axi_rmem15_ARREADY,
  m_axi_rmem15_ARSIZE,
  m_axi_rmem15_ARVALID,
  m_axi_rmem15_AWADDR,
  m_axi_rmem15_AWBURST,
  m_axi_rmem15_AWCACHE,
  m_axi_rmem15_AWID,
  m_axi_rmem15_AWLEN,
  m_axi_rmem15_AWLOCK,
  m_axi_rmem15_AWPROT,
  m_axi_rmem15_AWQOS,
  m_axi_rmem15_AWREADY,
  m_axi_rmem15_AWSIZE,
  m_axi_rmem15_AWVALID,
  m_axi_rmem15_BID,
  m_axi_rmem15_BREADY,
  m_axi_rmem15_BRESP,
  m_axi_rmem15_BVALID,
  m_axi_rmem15_RDATA,
  m_axi_rmem15_RID,
  m_axi_rmem15_RLAST,
  m_axi_rmem15_RREADY,
  m_axi_rmem15_RRESP,
  m_axi_rmem15_RVALID,
  m_axi_rmem15_WDATA,
  m_axi_rmem15_WLAST,
  m_axi_rmem15_WREADY,
  m_axi_rmem15_WSTRB,
  m_axi_rmem15_WVALID,
  m_axi_rmem16_ARADDR,
  m_axi_rmem16_ARBURST,
  m_axi_rmem16_ARCACHE,
  m_axi_rmem16_ARID,
  m_axi_rmem16_ARLEN,
  m_axi_rmem16_ARLOCK,
  m_axi_rmem16_ARPROT,
  m_axi_rmem16_ARQOS,
  m_axi_rmem16_ARREADY,
  m_axi_rmem16_ARSIZE,
  m_axi_rmem16_ARVALID,
  m_axi_rmem16_AWADDR,
  m_axi_rmem16_AWBURST,
  m_axi_rmem16_AWCACHE,
  m_axi_rmem16_AWID,
  m_axi_rmem16_AWLEN,
  m_axi_rmem16_AWLOCK,
  m_axi_rmem16_AWPROT,
  m_axi_rmem16_AWQOS,
  m_axi_rmem16_AWREADY,
  m_axi_rmem16_AWSIZE,
  m_axi_rmem16_AWVALID,
  m_axi_rmem16_BID,
  m_axi_rmem16_BREADY,
  m_axi_rmem16_BRESP,
  m_axi_rmem16_BVALID,
  m_axi_rmem16_RDATA,
  m_axi_rmem16_RID,
  m_axi_rmem16_RLAST,
  m_axi_rmem16_RREADY,
  m_axi_rmem16_RRESP,
  m_axi_rmem16_RVALID,
  m_axi_rmem16_WDATA,
  m_axi_rmem16_WLAST,
  m_axi_rmem16_WREADY,
  m_axi_rmem16_WSTRB,
  m_axi_rmem16_WVALID,
  m_axi_rmem17_ARADDR,
  m_axi_rmem17_ARBURST,
  m_axi_rmem17_ARCACHE,
  m_axi_rmem17_ARID,
  m_axi_rmem17_ARLEN,
  m_axi_rmem17_ARLOCK,
  m_axi_rmem17_ARPROT,
  m_axi_rmem17_ARQOS,
  m_axi_rmem17_ARREADY,
  m_axi_rmem17_ARSIZE,
  m_axi_rmem17_ARVALID,
  m_axi_rmem17_AWADDR,
  m_axi_rmem17_AWBURST,
  m_axi_rmem17_AWCACHE,
  m_axi_rmem17_AWID,
  m_axi_rmem17_AWLEN,
  m_axi_rmem17_AWLOCK,
  m_axi_rmem17_AWPROT,
  m_axi_rmem17_AWQOS,
  m_axi_rmem17_AWREADY,
  m_axi_rmem17_AWSIZE,
  m_axi_rmem17_AWVALID,
  m_axi_rmem17_BID,
  m_axi_rmem17_BREADY,
  m_axi_rmem17_BRESP,
  m_axi_rmem17_BVALID,
  m_axi_rmem17_RDATA,
  m_axi_rmem17_RID,
  m_axi_rmem17_RLAST,
  m_axi_rmem17_RREADY,
  m_axi_rmem17_RRESP,
  m_axi_rmem17_RVALID,
  m_axi_rmem17_WDATA,
  m_axi_rmem17_WLAST,
  m_axi_rmem17_WREADY,
  m_axi_rmem17_WSTRB,
  m_axi_rmem17_WVALID,
  m_axi_rmem18_ARADDR,
  m_axi_rmem18_ARBURST,
  m_axi_rmem18_ARCACHE,
  m_axi_rmem18_ARID,
  m_axi_rmem18_ARLEN,
  m_axi_rmem18_ARLOCK,
  m_axi_rmem18_ARPROT,
  m_axi_rmem18_ARQOS,
  m_axi_rmem18_ARREADY,
  m_axi_rmem18_ARSIZE,
  m_axi_rmem18_ARVALID,
  m_axi_rmem18_AWADDR,
  m_axi_rmem18_AWBURST,
  m_axi_rmem18_AWCACHE,
  m_axi_rmem18_AWID,
  m_axi_rmem18_AWLEN,
  m_axi_rmem18_AWLOCK,
  m_axi_rmem18_AWPROT,
  m_axi_rmem18_AWQOS,
  m_axi_rmem18_AWREADY,
  m_axi_rmem18_AWSIZE,
  m_axi_rmem18_AWVALID,
  m_axi_rmem18_BID,
  m_axi_rmem18_BREADY,
  m_axi_rmem18_BRESP,
  m_axi_rmem18_BVALID,
  m_axi_rmem18_RDATA,
  m_axi_rmem18_RID,
  m_axi_rmem18_RLAST,
  m_axi_rmem18_RREADY,
  m_axi_rmem18_RRESP,
  m_axi_rmem18_RVALID,
  m_axi_rmem18_WDATA,
  m_axi_rmem18_WLAST,
  m_axi_rmem18_WREADY,
  m_axi_rmem18_WSTRB,
  m_axi_rmem18_WVALID,
  m_axi_rmem19_ARADDR,
  m_axi_rmem19_ARBURST,
  m_axi_rmem19_ARCACHE,
  m_axi_rmem19_ARID,
  m_axi_rmem19_ARLEN,
  m_axi_rmem19_ARLOCK,
  m_axi_rmem19_ARPROT,
  m_axi_rmem19_ARQOS,
  m_axi_rmem19_ARREADY,
  m_axi_rmem19_ARSIZE,
  m_axi_rmem19_ARVALID,
  m_axi_rmem19_AWADDR,
  m_axi_rmem19_AWBURST,
  m_axi_rmem19_AWCACHE,
  m_axi_rmem19_AWID,
  m_axi_rmem19_AWLEN,
  m_axi_rmem19_AWLOCK,
  m_axi_rmem19_AWPROT,
  m_axi_rmem19_AWQOS,
  m_axi_rmem19_AWREADY,
  m_axi_rmem19_AWSIZE,
  m_axi_rmem19_AWVALID,
  m_axi_rmem19_BID,
  m_axi_rmem19_BREADY,
  m_axi_rmem19_BRESP,
  m_axi_rmem19_BVALID,
  m_axi_rmem19_RDATA,
  m_axi_rmem19_RID,
  m_axi_rmem19_RLAST,
  m_axi_rmem19_RREADY,
  m_axi_rmem19_RRESP,
  m_axi_rmem19_RVALID,
  m_axi_rmem19_WDATA,
  m_axi_rmem19_WLAST,
  m_axi_rmem19_WREADY,
  m_axi_rmem19_WSTRB,
  m_axi_rmem19_WVALID,
  m_axi_rmem20_ARADDR,
  m_axi_rmem20_ARBURST,
  m_axi_rmem20_ARCACHE,
  m_axi_rmem20_ARID,
  m_axi_rmem20_ARLEN,
  m_axi_rmem20_ARLOCK,
  m_axi_rmem20_ARPROT,
  m_axi_rmem20_ARQOS,
  m_axi_rmem20_ARREADY,
  m_axi_rmem20_ARSIZE,
  m_axi_rmem20_ARVALID,
  m_axi_rmem20_AWADDR,
  m_axi_rmem20_AWBURST,
  m_axi_rmem20_AWCACHE,
  m_axi_rmem20_AWID,
  m_axi_rmem20_AWLEN,
  m_axi_rmem20_AWLOCK,
  m_axi_rmem20_AWPROT,
  m_axi_rmem20_AWQOS,
  m_axi_rmem20_AWREADY,
  m_axi_rmem20_AWSIZE,
  m_axi_rmem20_AWVALID,
  m_axi_rmem20_BID,
  m_axi_rmem20_BREADY,
  m_axi_rmem20_BRESP,
  m_axi_rmem20_BVALID,
  m_axi_rmem20_RDATA,
  m_axi_rmem20_RID,
  m_axi_rmem20_RLAST,
  m_axi_rmem20_RREADY,
  m_axi_rmem20_RRESP,
  m_axi_rmem20_RVALID,
  m_axi_rmem20_WDATA,
  m_axi_rmem20_WLAST,
  m_axi_rmem20_WREADY,
  m_axi_rmem20_WSTRB,
  m_axi_rmem20_WVALID,
  m_axi_rmem21_ARADDR,
  m_axi_rmem21_ARBURST,
  m_axi_rmem21_ARCACHE,
  m_axi_rmem21_ARID,
  m_axi_rmem21_ARLEN,
  m_axi_rmem21_ARLOCK,
  m_axi_rmem21_ARPROT,
  m_axi_rmem21_ARQOS,
  m_axi_rmem21_ARREADY,
  m_axi_rmem21_ARSIZE,
  m_axi_rmem21_ARVALID,
  m_axi_rmem21_AWADDR,
  m_axi_rmem21_AWBURST,
  m_axi_rmem21_AWCACHE,
  m_axi_rmem21_AWID,
  m_axi_rmem21_AWLEN,
  m_axi_rmem21_AWLOCK,
  m_axi_rmem21_AWPROT,
  m_axi_rmem21_AWQOS,
  m_axi_rmem21_AWREADY,
  m_axi_rmem21_AWSIZE,
  m_axi_rmem21_AWVALID,
  m_axi_rmem21_BID,
  m_axi_rmem21_BREADY,
  m_axi_rmem21_BRESP,
  m_axi_rmem21_BVALID,
  m_axi_rmem21_RDATA,
  m_axi_rmem21_RID,
  m_axi_rmem21_RLAST,
  m_axi_rmem21_RREADY,
  m_axi_rmem21_RRESP,
  m_axi_rmem21_RVALID,
  m_axi_rmem21_WDATA,
  m_axi_rmem21_WLAST,
  m_axi_rmem21_WREADY,
  m_axi_rmem21_WSTRB,
  m_axi_rmem21_WVALID,
  m_axi_rmem22_ARADDR,
  m_axi_rmem22_ARBURST,
  m_axi_rmem22_ARCACHE,
  m_axi_rmem22_ARID,
  m_axi_rmem22_ARLEN,
  m_axi_rmem22_ARLOCK,
  m_axi_rmem22_ARPROT,
  m_axi_rmem22_ARQOS,
  m_axi_rmem22_ARREADY,
  m_axi_rmem22_ARSIZE,
  m_axi_rmem22_ARVALID,
  m_axi_rmem22_AWADDR,
  m_axi_rmem22_AWBURST,
  m_axi_rmem22_AWCACHE,
  m_axi_rmem22_AWID,
  m_axi_rmem22_AWLEN,
  m_axi_rmem22_AWLOCK,
  m_axi_rmem22_AWPROT,
  m_axi_rmem22_AWQOS,
  m_axi_rmem22_AWREADY,
  m_axi_rmem22_AWSIZE,
  m_axi_rmem22_AWVALID,
  m_axi_rmem22_BID,
  m_axi_rmem22_BREADY,
  m_axi_rmem22_BRESP,
  m_axi_rmem22_BVALID,
  m_axi_rmem22_RDATA,
  m_axi_rmem22_RID,
  m_axi_rmem22_RLAST,
  m_axi_rmem22_RREADY,
  m_axi_rmem22_RRESP,
  m_axi_rmem22_RVALID,
  m_axi_rmem22_WDATA,
  m_axi_rmem22_WLAST,
  m_axi_rmem22_WREADY,
  m_axi_rmem22_WSTRB,
  m_axi_rmem22_WVALID,
  m_axi_rmem23_ARADDR,
  m_axi_rmem23_ARBURST,
  m_axi_rmem23_ARCACHE,
  m_axi_rmem23_ARID,
  m_axi_rmem23_ARLEN,
  m_axi_rmem23_ARLOCK,
  m_axi_rmem23_ARPROT,
  m_axi_rmem23_ARQOS,
  m_axi_rmem23_ARREADY,
  m_axi_rmem23_ARSIZE,
  m_axi_rmem23_ARVALID,
  m_axi_rmem23_AWADDR,
  m_axi_rmem23_AWBURST,
  m_axi_rmem23_AWCACHE,
  m_axi_rmem23_AWID,
  m_axi_rmem23_AWLEN,
  m_axi_rmem23_AWLOCK,
  m_axi_rmem23_AWPROT,
  m_axi_rmem23_AWQOS,
  m_axi_rmem23_AWREADY,
  m_axi_rmem23_AWSIZE,
  m_axi_rmem23_AWVALID,
  m_axi_rmem23_BID,
  m_axi_rmem23_BREADY,
  m_axi_rmem23_BRESP,
  m_axi_rmem23_BVALID,
  m_axi_rmem23_RDATA,
  m_axi_rmem23_RID,
  m_axi_rmem23_RLAST,
  m_axi_rmem23_RREADY,
  m_axi_rmem23_RRESP,
  m_axi_rmem23_RVALID,
  m_axi_rmem23_WDATA,
  m_axi_rmem23_WLAST,
  m_axi_rmem23_WREADY,
  m_axi_rmem23_WSTRB,
  m_axi_rmem23_WVALID,
  m_axi_rmem24_ARADDR,
  m_axi_rmem24_ARBURST,
  m_axi_rmem24_ARCACHE,
  m_axi_rmem24_ARID,
  m_axi_rmem24_ARLEN,
  m_axi_rmem24_ARLOCK,
  m_axi_rmem24_ARPROT,
  m_axi_rmem24_ARQOS,
  m_axi_rmem24_ARREADY,
  m_axi_rmem24_ARSIZE,
  m_axi_rmem24_ARVALID,
  m_axi_rmem24_AWADDR,
  m_axi_rmem24_AWBURST,
  m_axi_rmem24_AWCACHE,
  m_axi_rmem24_AWID,
  m_axi_rmem24_AWLEN,
  m_axi_rmem24_AWLOCK,
  m_axi_rmem24_AWPROT,
  m_axi_rmem24_AWQOS,
  m_axi_rmem24_AWREADY,
  m_axi_rmem24_AWSIZE,
  m_axi_rmem24_AWVALID,
  m_axi_rmem24_BID,
  m_axi_rmem24_BREADY,
  m_axi_rmem24_BRESP,
  m_axi_rmem24_BVALID,
  m_axi_rmem24_RDATA,
  m_axi_rmem24_RID,
  m_axi_rmem24_RLAST,
  m_axi_rmem24_RREADY,
  m_axi_rmem24_RRESP,
  m_axi_rmem24_RVALID,
  m_axi_rmem24_WDATA,
  m_axi_rmem24_WLAST,
  m_axi_rmem24_WREADY,
  m_axi_rmem24_WSTRB,
  m_axi_rmem24_WVALID,
  m_axi_rmem25_ARADDR,
  m_axi_rmem25_ARBURST,
  m_axi_rmem25_ARCACHE,
  m_axi_rmem25_ARID,
  m_axi_rmem25_ARLEN,
  m_axi_rmem25_ARLOCK,
  m_axi_rmem25_ARPROT,
  m_axi_rmem25_ARQOS,
  m_axi_rmem25_ARREADY,
  m_axi_rmem25_ARSIZE,
  m_axi_rmem25_ARVALID,
  m_axi_rmem25_AWADDR,
  m_axi_rmem25_AWBURST,
  m_axi_rmem25_AWCACHE,
  m_axi_rmem25_AWID,
  m_axi_rmem25_AWLEN,
  m_axi_rmem25_AWLOCK,
  m_axi_rmem25_AWPROT,
  m_axi_rmem25_AWQOS,
  m_axi_rmem25_AWREADY,
  m_axi_rmem25_AWSIZE,
  m_axi_rmem25_AWVALID,
  m_axi_rmem25_BID,
  m_axi_rmem25_BREADY,
  m_axi_rmem25_BRESP,
  m_axi_rmem25_BVALID,
  m_axi_rmem25_RDATA,
  m_axi_rmem25_RID,
  m_axi_rmem25_RLAST,
  m_axi_rmem25_RREADY,
  m_axi_rmem25_RRESP,
  m_axi_rmem25_RVALID,
  m_axi_rmem25_WDATA,
  m_axi_rmem25_WLAST,
  m_axi_rmem25_WREADY,
  m_axi_rmem25_WSTRB,
  m_axi_rmem25_WVALID,
  m_axi_rmem26_ARADDR,
  m_axi_rmem26_ARBURST,
  m_axi_rmem26_ARCACHE,
  m_axi_rmem26_ARID,
  m_axi_rmem26_ARLEN,
  m_axi_rmem26_ARLOCK,
  m_axi_rmem26_ARPROT,
  m_axi_rmem26_ARQOS,
  m_axi_rmem26_ARREADY,
  m_axi_rmem26_ARSIZE,
  m_axi_rmem26_ARVALID,
  m_axi_rmem26_AWADDR,
  m_axi_rmem26_AWBURST,
  m_axi_rmem26_AWCACHE,
  m_axi_rmem26_AWID,
  m_axi_rmem26_AWLEN,
  m_axi_rmem26_AWLOCK,
  m_axi_rmem26_AWPROT,
  m_axi_rmem26_AWQOS,
  m_axi_rmem26_AWREADY,
  m_axi_rmem26_AWSIZE,
  m_axi_rmem26_AWVALID,
  m_axi_rmem26_BID,
  m_axi_rmem26_BREADY,
  m_axi_rmem26_BRESP,
  m_axi_rmem26_BVALID,
  m_axi_rmem26_RDATA,
  m_axi_rmem26_RID,
  m_axi_rmem26_RLAST,
  m_axi_rmem26_RREADY,
  m_axi_rmem26_RRESP,
  m_axi_rmem26_RVALID,
  m_axi_rmem26_WDATA,
  m_axi_rmem26_WLAST,
  m_axi_rmem26_WREADY,
  m_axi_rmem26_WSTRB,
  m_axi_rmem26_WVALID,
  m_axi_rmem27_ARADDR,
  m_axi_rmem27_ARBURST,
  m_axi_rmem27_ARCACHE,
  m_axi_rmem27_ARID,
  m_axi_rmem27_ARLEN,
  m_axi_rmem27_ARLOCK,
  m_axi_rmem27_ARPROT,
  m_axi_rmem27_ARQOS,
  m_axi_rmem27_ARREADY,
  m_axi_rmem27_ARSIZE,
  m_axi_rmem27_ARVALID,
  m_axi_rmem27_AWADDR,
  m_axi_rmem27_AWBURST,
  m_axi_rmem27_AWCACHE,
  m_axi_rmem27_AWID,
  m_axi_rmem27_AWLEN,
  m_axi_rmem27_AWLOCK,
  m_axi_rmem27_AWPROT,
  m_axi_rmem27_AWQOS,
  m_axi_rmem27_AWREADY,
  m_axi_rmem27_AWSIZE,
  m_axi_rmem27_AWVALID,
  m_axi_rmem27_BID,
  m_axi_rmem27_BREADY,
  m_axi_rmem27_BRESP,
  m_axi_rmem27_BVALID,
  m_axi_rmem27_RDATA,
  m_axi_rmem27_RID,
  m_axi_rmem27_RLAST,
  m_axi_rmem27_RREADY,
  m_axi_rmem27_RRESP,
  m_axi_rmem27_RVALID,
  m_axi_rmem27_WDATA,
  m_axi_rmem27_WLAST,
  m_axi_rmem27_WREADY,
  m_axi_rmem27_WSTRB,
  m_axi_rmem27_WVALID
);

  parameter C_S_AXI_CONTROL_DATA_WIDTH = 32;
  parameter C_S_AXI_CONTROL_ADDR_WIDTH = 9;
  parameter C_S_AXI_DATA_WIDTH = 32;
  parameter C_S_AXI_CONTROL_WSTRB_WIDTH = 32 / 8;
  parameter C_S_AXI_WSTRB_WIDTH = 32 / 8;
  (* RS_HS = "s_axi_control_AW.valid" *)input s_axi_control_AWVALID;
  (* RS_HS = "s_axi_control_AW.ready" *)output s_axi_control_AWREADY;
  (* RS_HS = "s_axi_control_AW.data" *)input [C_S_AXI_CONTROL_ADDR_WIDTH-1:0] s_axi_control_AWADDR;
  (* RS_HS = "s_axi_control_W.valid" *)input s_axi_control_WVALID;
  (* RS_HS = "s_axi_control_W.ready" *)output s_axi_control_WREADY;
  (* RS_HS = "s_axi_control_W.data" *)input [C_S_AXI_CONTROL_DATA_WIDTH-1:0] s_axi_control_WDATA;
  (* RS_HS = "s_axi_control_W.data" *)input [C_S_AXI_CONTROL_WSTRB_WIDTH-1:0] s_axi_control_WSTRB;
  (* RS_HS = "s_axi_control_AR.valid" *)input s_axi_control_ARVALID;
  (* RS_HS = "s_axi_control_AR.ready" *)output s_axi_control_ARREADY;
  (* RS_HS = "s_axi_control_AR.data" *)input [C_S_AXI_CONTROL_ADDR_WIDTH-1:0] s_axi_control_ARADDR;
  (* RS_HS = "s_axi_control_R.valid" *)output s_axi_control_RVALID;
  (* RS_HS = "s_axi_control_R.ready" *)input s_axi_control_RREADY;
  (* RS_HS = "s_axi_control_R.data" *)output [C_S_AXI_CONTROL_DATA_WIDTH-1:0] s_axi_control_RDATA;
  (* RS_HS = "s_axi_control_R.data" *)output [1:0] s_axi_control_RRESP;
  (* RS_HS = "s_axi_control_B.valid" *)output s_axi_control_BVALID;
  (* RS_HS = "s_axi_control_B.ready" *)input s_axi_control_BREADY;
  (* RS_HS = "s_axi_control_B.data" *)output [1:0] s_axi_control_BRESP;
  (* RS_CLK *)input ap_clk;
  (* RS_RST = "ff" *)input ap_rst_n;
  (* RS_FF = "interrupt" *)output interrupt;
  (* RS_HS = "m_axi_rmem0_AR.data" *)output [63:0] m_axi_rmem0_ARADDR;
  (* RS_HS = "m_axi_rmem0_AR.data" *)output [1:0] m_axi_rmem0_ARBURST;
  (* RS_HS = "m_axi_rmem0_AR.data" *)output [3:0] m_axi_rmem0_ARCACHE;
  (* RS_HS = "m_axi_rmem0_AR.data" *)output [1:0] m_axi_rmem0_ARID;
  (* RS_HS = "m_axi_rmem0_AR.data" *)output [7:0] m_axi_rmem0_ARLEN;
  (* RS_HS = "m_axi_rmem0_AR.data" *)output m_axi_rmem0_ARLOCK;
  (* RS_HS = "m_axi_rmem0_AR.data" *)output [2:0] m_axi_rmem0_ARPROT;
  (* RS_HS = "m_axi_rmem0_AR.data" *)output [3:0] m_axi_rmem0_ARQOS;
  (* RS_HS = "m_axi_rmem0_AR.ready" *)input m_axi_rmem0_ARREADY;
  (* RS_HS = "m_axi_rmem0_AR.data" *)output [2:0] m_axi_rmem0_ARSIZE;
  (* RS_HS = "m_axi_rmem0_AR.valid" *)output m_axi_rmem0_ARVALID;
  (* RS_HS = "m_axi_rmem0_AW.data" *)output [63:0] m_axi_rmem0_AWADDR;
  (* RS_HS = "m_axi_rmem0_AW.data" *)output [1:0] m_axi_rmem0_AWBURST;
  (* RS_HS = "m_axi_rmem0_AW.data" *)output [3:0] m_axi_rmem0_AWCACHE;
  (* RS_HS = "m_axi_rmem0_AW.data" *)output [1:0] m_axi_rmem0_AWID;
  (* RS_HS = "m_axi_rmem0_AW.data" *)output [7:0] m_axi_rmem0_AWLEN;
  (* RS_HS = "m_axi_rmem0_AW.data" *)output m_axi_rmem0_AWLOCK;
  (* RS_HS = "m_axi_rmem0_AW.data" *)output [2:0] m_axi_rmem0_AWPROT;
  (* RS_HS = "m_axi_rmem0_AW.data" *)output [3:0] m_axi_rmem0_AWQOS;
  (* RS_HS = "m_axi_rmem0_AW.ready" *)input m_axi_rmem0_AWREADY;
  (* RS_HS = "m_axi_rmem0_AW.data" *)output [2:0] m_axi_rmem0_AWSIZE;
  (* RS_HS = "m_axi_rmem0_AW.valid" *)output m_axi_rmem0_AWVALID;
  (* RS_HS = "m_axi_rmem0_B.data" *)input [1:0] m_axi_rmem0_BID;
  (* RS_HS = "m_axi_rmem0_B.ready" *)output m_axi_rmem0_BREADY;
  (* RS_HS = "m_axi_rmem0_B.data" *)input [1:0] m_axi_rmem0_BRESP;
  (* RS_HS = "m_axi_rmem0_B.valid" *)input m_axi_rmem0_BVALID;
  (* RS_HS = "m_axi_rmem0_R.data" *)input [511:0] m_axi_rmem0_RDATA;
  (* RS_HS = "m_axi_rmem0_R.data" *)input [1:0] m_axi_rmem0_RID;
  (* RS_HS = "m_axi_rmem0_R.data" *)input m_axi_rmem0_RLAST;
  (* RS_HS = "m_axi_rmem0_R.ready" *)output m_axi_rmem0_RREADY;
  (* RS_HS = "m_axi_rmem0_R.data" *)input [1:0] m_axi_rmem0_RRESP;
  (* RS_HS = "m_axi_rmem0_R.valid" *)input m_axi_rmem0_RVALID;
  (* RS_HS = "m_axi_rmem0_W.data" *)output [511:0] m_axi_rmem0_WDATA;
  (* RS_HS = "m_axi_rmem0_W.data" *)output m_axi_rmem0_WLAST;
  (* RS_HS = "m_axi_rmem0_W.ready" *)input m_axi_rmem0_WREADY;
  (* RS_HS = "m_axi_rmem0_W.data" *)output [63:0] m_axi_rmem0_WSTRB;
  (* RS_HS = "m_axi_rmem0_W.valid" *)output m_axi_rmem0_WVALID;
  (* RS_HS = "m_axi_rmem1_AR.data" *)output [63:0] m_axi_rmem1_ARADDR;
  (* RS_HS = "m_axi_rmem1_AR.data" *)output [1:0] m_axi_rmem1_ARBURST;
  (* RS_HS = "m_axi_rmem1_AR.data" *)output [3:0] m_axi_rmem1_ARCACHE;
  (* RS_HS = "m_axi_rmem1_AR.data" *)output [1:0] m_axi_rmem1_ARID;
  (* RS_HS = "m_axi_rmem1_AR.data" *)output [7:0] m_axi_rmem1_ARLEN;
  (* RS_HS = "m_axi_rmem1_AR.data" *)output m_axi_rmem1_ARLOCK;
  (* RS_HS = "m_axi_rmem1_AR.data" *)output [2:0] m_axi_rmem1_ARPROT;
  (* RS_HS = "m_axi_rmem1_AR.data" *)output [3:0] m_axi_rmem1_ARQOS;
  (* RS_HS = "m_axi_rmem1_AR.ready" *)input m_axi_rmem1_ARREADY;
  (* RS_HS = "m_axi_rmem1_AR.data" *)output [2:0] m_axi_rmem1_ARSIZE;
  (* RS_HS = "m_axi_rmem1_AR.valid" *)output m_axi_rmem1_ARVALID;
  (* RS_HS = "m_axi_rmem1_AW.data" *)output [63:0] m_axi_rmem1_AWADDR;
  (* RS_HS = "m_axi_rmem1_AW.data" *)output [1:0] m_axi_rmem1_AWBURST;
  (* RS_HS = "m_axi_rmem1_AW.data" *)output [3:0] m_axi_rmem1_AWCACHE;
  (* RS_HS = "m_axi_rmem1_AW.data" *)output [1:0] m_axi_rmem1_AWID;
  (* RS_HS = "m_axi_rmem1_AW.data" *)output [7:0] m_axi_rmem1_AWLEN;
  (* RS_HS = "m_axi_rmem1_AW.data" *)output m_axi_rmem1_AWLOCK;
  (* RS_HS = "m_axi_rmem1_AW.data" *)output [2:0] m_axi_rmem1_AWPROT;
  (* RS_HS = "m_axi_rmem1_AW.data" *)output [3:0] m_axi_rmem1_AWQOS;
  (* RS_HS = "m_axi_rmem1_AW.ready" *)input m_axi_rmem1_AWREADY;
  (* RS_HS = "m_axi_rmem1_AW.data" *)output [2:0] m_axi_rmem1_AWSIZE;
  (* RS_HS = "m_axi_rmem1_AW.valid" *)output m_axi_rmem1_AWVALID;
  (* RS_HS = "m_axi_rmem1_B.data" *)input [1:0] m_axi_rmem1_BID;
  (* RS_HS = "m_axi_rmem1_B.ready" *)output m_axi_rmem1_BREADY;
  (* RS_HS = "m_axi_rmem1_B.data" *)input [1:0] m_axi_rmem1_BRESP;
  (* RS_HS = "m_axi_rmem1_B.valid" *)input m_axi_rmem1_BVALID;
  (* RS_HS = "m_axi_rmem1_R.data" *)input [511:0] m_axi_rmem1_RDATA;
  (* RS_HS = "m_axi_rmem1_R.data" *)input [1:0] m_axi_rmem1_RID;
  (* RS_HS = "m_axi_rmem1_R.data" *)input m_axi_rmem1_RLAST;
  (* RS_HS = "m_axi_rmem1_R.ready" *)output m_axi_rmem1_RREADY;
  (* RS_HS = "m_axi_rmem1_R.data" *)input [1:0] m_axi_rmem1_RRESP;
  (* RS_HS = "m_axi_rmem1_R.valid" *)input m_axi_rmem1_RVALID;
  (* RS_HS = "m_axi_rmem1_W.data" *)output [511:0] m_axi_rmem1_WDATA;
  (* RS_HS = "m_axi_rmem1_W.data" *)output m_axi_rmem1_WLAST;
  (* RS_HS = "m_axi_rmem1_W.ready" *)input m_axi_rmem1_WREADY;
  (* RS_HS = "m_axi_rmem1_W.data" *)output [63:0] m_axi_rmem1_WSTRB;
  (* RS_HS = "m_axi_rmem1_W.valid" *)output m_axi_rmem1_WVALID;
  (* RS_HS = "m_axi_rmem2_AR.data" *)output [63:0] m_axi_rmem2_ARADDR;
  (* RS_HS = "m_axi_rmem2_AR.data" *)output [1:0] m_axi_rmem2_ARBURST;
  (* RS_HS = "m_axi_rmem2_AR.data" *)output [3:0] m_axi_rmem2_ARCACHE;
  (* RS_HS = "m_axi_rmem2_AR.data" *)output [1:0] m_axi_rmem2_ARID;
  (* RS_HS = "m_axi_rmem2_AR.data" *)output [7:0] m_axi_rmem2_ARLEN;
  (* RS_HS = "m_axi_rmem2_AR.data" *)output m_axi_rmem2_ARLOCK;
  (* RS_HS = "m_axi_rmem2_AR.data" *)output [2:0] m_axi_rmem2_ARPROT;
  (* RS_HS = "m_axi_rmem2_AR.data" *)output [3:0] m_axi_rmem2_ARQOS;
  (* RS_HS = "m_axi_rmem2_AR.ready" *)input m_axi_rmem2_ARREADY;
  (* RS_HS = "m_axi_rmem2_AR.data" *)output [2:0] m_axi_rmem2_ARSIZE;
  (* RS_HS = "m_axi_rmem2_AR.valid" *)output m_axi_rmem2_ARVALID;
  (* RS_HS = "m_axi_rmem2_AW.data" *)output [63:0] m_axi_rmem2_AWADDR;
  (* RS_HS = "m_axi_rmem2_AW.data" *)output [1:0] m_axi_rmem2_AWBURST;
  (* RS_HS = "m_axi_rmem2_AW.data" *)output [3:0] m_axi_rmem2_AWCACHE;
  (* RS_HS = "m_axi_rmem2_AW.data" *)output [1:0] m_axi_rmem2_AWID;
  (* RS_HS = "m_axi_rmem2_AW.data" *)output [7:0] m_axi_rmem2_AWLEN;
  (* RS_HS = "m_axi_rmem2_AW.data" *)output m_axi_rmem2_AWLOCK;
  (* RS_HS = "m_axi_rmem2_AW.data" *)output [2:0] m_axi_rmem2_AWPROT;
  (* RS_HS = "m_axi_rmem2_AW.data" *)output [3:0] m_axi_rmem2_AWQOS;
  (* RS_HS = "m_axi_rmem2_AW.ready" *)input m_axi_rmem2_AWREADY;
  (* RS_HS = "m_axi_rmem2_AW.data" *)output [2:0] m_axi_rmem2_AWSIZE;
  (* RS_HS = "m_axi_rmem2_AW.valid" *)output m_axi_rmem2_AWVALID;
  (* RS_HS = "m_axi_rmem2_B.data" *)input [1:0] m_axi_rmem2_BID;
  (* RS_HS = "m_axi_rmem2_B.ready" *)output m_axi_rmem2_BREADY;
  (* RS_HS = "m_axi_rmem2_B.data" *)input [1:0] m_axi_rmem2_BRESP;
  (* RS_HS = "m_axi_rmem2_B.valid" *)input m_axi_rmem2_BVALID;
  (* RS_HS = "m_axi_rmem2_R.data" *)input [511:0] m_axi_rmem2_RDATA;
  (* RS_HS = "m_axi_rmem2_R.data" *)input [1:0] m_axi_rmem2_RID;
  (* RS_HS = "m_axi_rmem2_R.data" *)input m_axi_rmem2_RLAST;
  (* RS_HS = "m_axi_rmem2_R.ready" *)output m_axi_rmem2_RREADY;
  (* RS_HS = "m_axi_rmem2_R.data" *)input [1:0] m_axi_rmem2_RRESP;
  (* RS_HS = "m_axi_rmem2_R.valid" *)input m_axi_rmem2_RVALID;
  (* RS_HS = "m_axi_rmem2_W.data" *)output [511:0] m_axi_rmem2_WDATA;
  (* RS_HS = "m_axi_rmem2_W.data" *)output m_axi_rmem2_WLAST;
  (* RS_HS = "m_axi_rmem2_W.ready" *)input m_axi_rmem2_WREADY;
  (* RS_HS = "m_axi_rmem2_W.data" *)output [63:0] m_axi_rmem2_WSTRB;
  (* RS_HS = "m_axi_rmem2_W.valid" *)output m_axi_rmem2_WVALID;
  (* RS_HS = "m_axi_rmem3_AR.data" *)output [63:0] m_axi_rmem3_ARADDR;
  (* RS_HS = "m_axi_rmem3_AR.data" *)output [1:0] m_axi_rmem3_ARBURST;
  (* RS_HS = "m_axi_rmem3_AR.data" *)output [3:0] m_axi_rmem3_ARCACHE;
  (* RS_HS = "m_axi_rmem3_AR.data" *)output [1:0] m_axi_rmem3_ARID;
  (* RS_HS = "m_axi_rmem3_AR.data" *)output [7:0] m_axi_rmem3_ARLEN;
  (* RS_HS = "m_axi_rmem3_AR.data" *)output m_axi_rmem3_ARLOCK;
  (* RS_HS = "m_axi_rmem3_AR.data" *)output [2:0] m_axi_rmem3_ARPROT;
  (* RS_HS = "m_axi_rmem3_AR.data" *)output [3:0] m_axi_rmem3_ARQOS;
  (* RS_HS = "m_axi_rmem3_AR.ready" *)input m_axi_rmem3_ARREADY;
  (* RS_HS = "m_axi_rmem3_AR.data" *)output [2:0] m_axi_rmem3_ARSIZE;
  (* RS_HS = "m_axi_rmem3_AR.valid" *)output m_axi_rmem3_ARVALID;
  (* RS_HS = "m_axi_rmem3_AW.data" *)output [63:0] m_axi_rmem3_AWADDR;
  (* RS_HS = "m_axi_rmem3_AW.data" *)output [1:0] m_axi_rmem3_AWBURST;
  (* RS_HS = "m_axi_rmem3_AW.data" *)output [3:0] m_axi_rmem3_AWCACHE;
  (* RS_HS = "m_axi_rmem3_AW.data" *)output [1:0] m_axi_rmem3_AWID;
  (* RS_HS = "m_axi_rmem3_AW.data" *)output [7:0] m_axi_rmem3_AWLEN;
  (* RS_HS = "m_axi_rmem3_AW.data" *)output m_axi_rmem3_AWLOCK;
  (* RS_HS = "m_axi_rmem3_AW.data" *)output [2:0] m_axi_rmem3_AWPROT;
  (* RS_HS = "m_axi_rmem3_AW.data" *)output [3:0] m_axi_rmem3_AWQOS;
  (* RS_HS = "m_axi_rmem3_AW.ready" *)input m_axi_rmem3_AWREADY;
  (* RS_HS = "m_axi_rmem3_AW.data" *)output [2:0] m_axi_rmem3_AWSIZE;
  (* RS_HS = "m_axi_rmem3_AW.valid" *)output m_axi_rmem3_AWVALID;
  (* RS_HS = "m_axi_rmem3_B.data" *)input [1:0] m_axi_rmem3_BID;
  (* RS_HS = "m_axi_rmem3_B.ready" *)output m_axi_rmem3_BREADY;
  (* RS_HS = "m_axi_rmem3_B.data" *)input [1:0] m_axi_rmem3_BRESP;
  (* RS_HS = "m_axi_rmem3_B.valid" *)input m_axi_rmem3_BVALID;
  (* RS_HS = "m_axi_rmem3_R.data" *)input [511:0] m_axi_rmem3_RDATA;
  (* RS_HS = "m_axi_rmem3_R.data" *)input [1:0] m_axi_rmem3_RID;
  (* RS_HS = "m_axi_rmem3_R.data" *)input m_axi_rmem3_RLAST;
  (* RS_HS = "m_axi_rmem3_R.ready" *)output m_axi_rmem3_RREADY;
  (* RS_HS = "m_axi_rmem3_R.data" *)input [1:0] m_axi_rmem3_RRESP;
  (* RS_HS = "m_axi_rmem3_R.valid" *)input m_axi_rmem3_RVALID;
  (* RS_HS = "m_axi_rmem3_W.data" *)output [511:0] m_axi_rmem3_WDATA;
  (* RS_HS = "m_axi_rmem3_W.data" *)output m_axi_rmem3_WLAST;
  (* RS_HS = "m_axi_rmem3_W.ready" *)input m_axi_rmem3_WREADY;
  (* RS_HS = "m_axi_rmem3_W.data" *)output [63:0] m_axi_rmem3_WSTRB;
  (* RS_HS = "m_axi_rmem3_W.valid" *)output m_axi_rmem3_WVALID;
  (* RS_HS = "m_axi_rmem4_AR.data" *)output [63:0] m_axi_rmem4_ARADDR;
  (* RS_HS = "m_axi_rmem4_AR.data" *)output [1:0] m_axi_rmem4_ARBURST;
  (* RS_HS = "m_axi_rmem4_AR.data" *)output [3:0] m_axi_rmem4_ARCACHE;
  (* RS_HS = "m_axi_rmem4_AR.data" *)output [1:0] m_axi_rmem4_ARID;
  (* RS_HS = "m_axi_rmem4_AR.data" *)output [7:0] m_axi_rmem4_ARLEN;
  (* RS_HS = "m_axi_rmem4_AR.data" *)output m_axi_rmem4_ARLOCK;
  (* RS_HS = "m_axi_rmem4_AR.data" *)output [2:0] m_axi_rmem4_ARPROT;
  (* RS_HS = "m_axi_rmem4_AR.data" *)output [3:0] m_axi_rmem4_ARQOS;
  (* RS_HS = "m_axi_rmem4_AR.ready" *)input m_axi_rmem4_ARREADY;
  (* RS_HS = "m_axi_rmem4_AR.data" *)output [2:0] m_axi_rmem4_ARSIZE;
  (* RS_HS = "m_axi_rmem4_AR.valid" *)output m_axi_rmem4_ARVALID;
  (* RS_HS = "m_axi_rmem4_AW.data" *)output [63:0] m_axi_rmem4_AWADDR;
  (* RS_HS = "m_axi_rmem4_AW.data" *)output [1:0] m_axi_rmem4_AWBURST;
  (* RS_HS = "m_axi_rmem4_AW.data" *)output [3:0] m_axi_rmem4_AWCACHE;
  (* RS_HS = "m_axi_rmem4_AW.data" *)output [1:0] m_axi_rmem4_AWID;
  (* RS_HS = "m_axi_rmem4_AW.data" *)output [7:0] m_axi_rmem4_AWLEN;
  (* RS_HS = "m_axi_rmem4_AW.data" *)output m_axi_rmem4_AWLOCK;
  (* RS_HS = "m_axi_rmem4_AW.data" *)output [2:0] m_axi_rmem4_AWPROT;
  (* RS_HS = "m_axi_rmem4_AW.data" *)output [3:0] m_axi_rmem4_AWQOS;
  (* RS_HS = "m_axi_rmem4_AW.ready" *)input m_axi_rmem4_AWREADY;
  (* RS_HS = "m_axi_rmem4_AW.data" *)output [2:0] m_axi_rmem4_AWSIZE;
  (* RS_HS = "m_axi_rmem4_AW.valid" *)output m_axi_rmem4_AWVALID;
  (* RS_HS = "m_axi_rmem4_B.data" *)input [1:0] m_axi_rmem4_BID;
  (* RS_HS = "m_axi_rmem4_B.ready" *)output m_axi_rmem4_BREADY;
  (* RS_HS = "m_axi_rmem4_B.data" *)input [1:0] m_axi_rmem4_BRESP;
  (* RS_HS = "m_axi_rmem4_B.valid" *)input m_axi_rmem4_BVALID;
  (* RS_HS = "m_axi_rmem4_R.data" *)input [511:0] m_axi_rmem4_RDATA;
  (* RS_HS = "m_axi_rmem4_R.data" *)input [1:0] m_axi_rmem4_RID;
  (* RS_HS = "m_axi_rmem4_R.data" *)input m_axi_rmem4_RLAST;
  (* RS_HS = "m_axi_rmem4_R.ready" *)output m_axi_rmem4_RREADY;
  (* RS_HS = "m_axi_rmem4_R.data" *)input [1:0] m_axi_rmem4_RRESP;
  (* RS_HS = "m_axi_rmem4_R.valid" *)input m_axi_rmem4_RVALID;
  (* RS_HS = "m_axi_rmem4_W.data" *)output [511:0] m_axi_rmem4_WDATA;
  (* RS_HS = "m_axi_rmem4_W.data" *)output m_axi_rmem4_WLAST;
  (* RS_HS = "m_axi_rmem4_W.ready" *)input m_axi_rmem4_WREADY;
  (* RS_HS = "m_axi_rmem4_W.data" *)output [63:0] m_axi_rmem4_WSTRB;
  (* RS_HS = "m_axi_rmem4_W.valid" *)output m_axi_rmem4_WVALID;
  (* RS_HS = "m_axi_rmem5_AR.data" *)output [63:0] m_axi_rmem5_ARADDR;
  (* RS_HS = "m_axi_rmem5_AR.data" *)output [1:0] m_axi_rmem5_ARBURST;
  (* RS_HS = "m_axi_rmem5_AR.data" *)output [3:0] m_axi_rmem5_ARCACHE;
  (* RS_HS = "m_axi_rmem5_AR.data" *)output [1:0] m_axi_rmem5_ARID;
  (* RS_HS = "m_axi_rmem5_AR.data" *)output [7:0] m_axi_rmem5_ARLEN;
  (* RS_HS = "m_axi_rmem5_AR.data" *)output m_axi_rmem5_ARLOCK;
  (* RS_HS = "m_axi_rmem5_AR.data" *)output [2:0] m_axi_rmem5_ARPROT;
  (* RS_HS = "m_axi_rmem5_AR.data" *)output [3:0] m_axi_rmem5_ARQOS;
  (* RS_HS = "m_axi_rmem5_AR.ready" *)input m_axi_rmem5_ARREADY;
  (* RS_HS = "m_axi_rmem5_AR.data" *)output [2:0] m_axi_rmem5_ARSIZE;
  (* RS_HS = "m_axi_rmem5_AR.valid" *)output m_axi_rmem5_ARVALID;
  (* RS_HS = "m_axi_rmem5_AW.data" *)output [63:0] m_axi_rmem5_AWADDR;
  (* RS_HS = "m_axi_rmem5_AW.data" *)output [1:0] m_axi_rmem5_AWBURST;
  (* RS_HS = "m_axi_rmem5_AW.data" *)output [3:0] m_axi_rmem5_AWCACHE;
  (* RS_HS = "m_axi_rmem5_AW.data" *)output [1:0] m_axi_rmem5_AWID;
  (* RS_HS = "m_axi_rmem5_AW.data" *)output [7:0] m_axi_rmem5_AWLEN;
  (* RS_HS = "m_axi_rmem5_AW.data" *)output m_axi_rmem5_AWLOCK;
  (* RS_HS = "m_axi_rmem5_AW.data" *)output [2:0] m_axi_rmem5_AWPROT;
  (* RS_HS = "m_axi_rmem5_AW.data" *)output [3:0] m_axi_rmem5_AWQOS;
  (* RS_HS = "m_axi_rmem5_AW.ready" *)input m_axi_rmem5_AWREADY;
  (* RS_HS = "m_axi_rmem5_AW.data" *)output [2:0] m_axi_rmem5_AWSIZE;
  (* RS_HS = "m_axi_rmem5_AW.valid" *)output m_axi_rmem5_AWVALID;
  (* RS_HS = "m_axi_rmem5_B.data" *)input [1:0] m_axi_rmem5_BID;
  (* RS_HS = "m_axi_rmem5_B.ready" *)output m_axi_rmem5_BREADY;
  (* RS_HS = "m_axi_rmem5_B.data" *)input [1:0] m_axi_rmem5_BRESP;
  (* RS_HS = "m_axi_rmem5_B.valid" *)input m_axi_rmem5_BVALID;
  (* RS_HS = "m_axi_rmem5_R.data" *)input [511:0] m_axi_rmem5_RDATA;
  (* RS_HS = "m_axi_rmem5_R.data" *)input [1:0] m_axi_rmem5_RID;
  (* RS_HS = "m_axi_rmem5_R.data" *)input m_axi_rmem5_RLAST;
  (* RS_HS = "m_axi_rmem5_R.ready" *)output m_axi_rmem5_RREADY;
  (* RS_HS = "m_axi_rmem5_R.data" *)input [1:0] m_axi_rmem5_RRESP;
  (* RS_HS = "m_axi_rmem5_R.valid" *)input m_axi_rmem5_RVALID;
  (* RS_HS = "m_axi_rmem5_W.data" *)output [511:0] m_axi_rmem5_WDATA;
  (* RS_HS = "m_axi_rmem5_W.data" *)output m_axi_rmem5_WLAST;
  (* RS_HS = "m_axi_rmem5_W.ready" *)input m_axi_rmem5_WREADY;
  (* RS_HS = "m_axi_rmem5_W.data" *)output [63:0] m_axi_rmem5_WSTRB;
  (* RS_HS = "m_axi_rmem5_W.valid" *)output m_axi_rmem5_WVALID;
  (* RS_HS = "m_axi_rmem6_AR.data" *)output [63:0] m_axi_rmem6_ARADDR;
  (* RS_HS = "m_axi_rmem6_AR.data" *)output [1:0] m_axi_rmem6_ARBURST;
  (* RS_HS = "m_axi_rmem6_AR.data" *)output [3:0] m_axi_rmem6_ARCACHE;
  (* RS_HS = "m_axi_rmem6_AR.data" *)output [1:0] m_axi_rmem6_ARID;
  (* RS_HS = "m_axi_rmem6_AR.data" *)output [7:0] m_axi_rmem6_ARLEN;
  (* RS_HS = "m_axi_rmem6_AR.data" *)output m_axi_rmem6_ARLOCK;
  (* RS_HS = "m_axi_rmem6_AR.data" *)output [2:0] m_axi_rmem6_ARPROT;
  (* RS_HS = "m_axi_rmem6_AR.data" *)output [3:0] m_axi_rmem6_ARQOS;
  (* RS_HS = "m_axi_rmem6_AR.ready" *)input m_axi_rmem6_ARREADY;
  (* RS_HS = "m_axi_rmem6_AR.data" *)output [2:0] m_axi_rmem6_ARSIZE;
  (* RS_HS = "m_axi_rmem6_AR.valid" *)output m_axi_rmem6_ARVALID;
  (* RS_HS = "m_axi_rmem6_AW.data" *)output [63:0] m_axi_rmem6_AWADDR;
  (* RS_HS = "m_axi_rmem6_AW.data" *)output [1:0] m_axi_rmem6_AWBURST;
  (* RS_HS = "m_axi_rmem6_AW.data" *)output [3:0] m_axi_rmem6_AWCACHE;
  (* RS_HS = "m_axi_rmem6_AW.data" *)output [1:0] m_axi_rmem6_AWID;
  (* RS_HS = "m_axi_rmem6_AW.data" *)output [7:0] m_axi_rmem6_AWLEN;
  (* RS_HS = "m_axi_rmem6_AW.data" *)output m_axi_rmem6_AWLOCK;
  (* RS_HS = "m_axi_rmem6_AW.data" *)output [2:0] m_axi_rmem6_AWPROT;
  (* RS_HS = "m_axi_rmem6_AW.data" *)output [3:0] m_axi_rmem6_AWQOS;
  (* RS_HS = "m_axi_rmem6_AW.ready" *)input m_axi_rmem6_AWREADY;
  (* RS_HS = "m_axi_rmem6_AW.data" *)output [2:0] m_axi_rmem6_AWSIZE;
  (* RS_HS = "m_axi_rmem6_AW.valid" *)output m_axi_rmem6_AWVALID;
  (* RS_HS = "m_axi_rmem6_B.data" *)input [1:0] m_axi_rmem6_BID;
  (* RS_HS = "m_axi_rmem6_B.ready" *)output m_axi_rmem6_BREADY;
  (* RS_HS = "m_axi_rmem6_B.data" *)input [1:0] m_axi_rmem6_BRESP;
  (* RS_HS = "m_axi_rmem6_B.valid" *)input m_axi_rmem6_BVALID;
  (* RS_HS = "m_axi_rmem6_R.data" *)input [511:0] m_axi_rmem6_RDATA;
  (* RS_HS = "m_axi_rmem6_R.data" *)input [1:0] m_axi_rmem6_RID;
  (* RS_HS = "m_axi_rmem6_R.data" *)input m_axi_rmem6_RLAST;
  (* RS_HS = "m_axi_rmem6_R.ready" *)output m_axi_rmem6_RREADY;
  (* RS_HS = "m_axi_rmem6_R.data" *)input [1:0] m_axi_rmem6_RRESP;
  (* RS_HS = "m_axi_rmem6_R.valid" *)input m_axi_rmem6_RVALID;
  (* RS_HS = "m_axi_rmem6_W.data" *)output [511:0] m_axi_rmem6_WDATA;
  (* RS_HS = "m_axi_rmem6_W.data" *)output m_axi_rmem6_WLAST;
  (* RS_HS = "m_axi_rmem6_W.ready" *)input m_axi_rmem6_WREADY;
  (* RS_HS = "m_axi_rmem6_W.data" *)output [63:0] m_axi_rmem6_WSTRB;
  (* RS_HS = "m_axi_rmem6_W.valid" *)output m_axi_rmem6_WVALID;
  (* RS_HS = "m_axi_rmem7_AR.data" *)output [63:0] m_axi_rmem7_ARADDR;
  (* RS_HS = "m_axi_rmem7_AR.data" *)output [1:0] m_axi_rmem7_ARBURST;
  (* RS_HS = "m_axi_rmem7_AR.data" *)output [3:0] m_axi_rmem7_ARCACHE;
  (* RS_HS = "m_axi_rmem7_AR.data" *)output [1:0] m_axi_rmem7_ARID;
  (* RS_HS = "m_axi_rmem7_AR.data" *)output [7:0] m_axi_rmem7_ARLEN;
  (* RS_HS = "m_axi_rmem7_AR.data" *)output m_axi_rmem7_ARLOCK;
  (* RS_HS = "m_axi_rmem7_AR.data" *)output [2:0] m_axi_rmem7_ARPROT;
  (* RS_HS = "m_axi_rmem7_AR.data" *)output [3:0] m_axi_rmem7_ARQOS;
  (* RS_HS = "m_axi_rmem7_AR.ready" *)input m_axi_rmem7_ARREADY;
  (* RS_HS = "m_axi_rmem7_AR.data" *)output [2:0] m_axi_rmem7_ARSIZE;
  (* RS_HS = "m_axi_rmem7_AR.valid" *)output m_axi_rmem7_ARVALID;
  (* RS_HS = "m_axi_rmem7_AW.data" *)output [63:0] m_axi_rmem7_AWADDR;
  (* RS_HS = "m_axi_rmem7_AW.data" *)output [1:0] m_axi_rmem7_AWBURST;
  (* RS_HS = "m_axi_rmem7_AW.data" *)output [3:0] m_axi_rmem7_AWCACHE;
  (* RS_HS = "m_axi_rmem7_AW.data" *)output [1:0] m_axi_rmem7_AWID;
  (* RS_HS = "m_axi_rmem7_AW.data" *)output [7:0] m_axi_rmem7_AWLEN;
  (* RS_HS = "m_axi_rmem7_AW.data" *)output m_axi_rmem7_AWLOCK;
  (* RS_HS = "m_axi_rmem7_AW.data" *)output [2:0] m_axi_rmem7_AWPROT;
  (* RS_HS = "m_axi_rmem7_AW.data" *)output [3:0] m_axi_rmem7_AWQOS;
  (* RS_HS = "m_axi_rmem7_AW.ready" *)input m_axi_rmem7_AWREADY;
  (* RS_HS = "m_axi_rmem7_AW.data" *)output [2:0] m_axi_rmem7_AWSIZE;
  (* RS_HS = "m_axi_rmem7_AW.valid" *)output m_axi_rmem7_AWVALID;
  (* RS_HS = "m_axi_rmem7_B.data" *)input [1:0] m_axi_rmem7_BID;
  (* RS_HS = "m_axi_rmem7_B.ready" *)output m_axi_rmem7_BREADY;
  (* RS_HS = "m_axi_rmem7_B.data" *)input [1:0] m_axi_rmem7_BRESP;
  (* RS_HS = "m_axi_rmem7_B.valid" *)input m_axi_rmem7_BVALID;
  (* RS_HS = "m_axi_rmem7_R.data" *)input [511:0] m_axi_rmem7_RDATA;
  (* RS_HS = "m_axi_rmem7_R.data" *)input [1:0] m_axi_rmem7_RID;
  (* RS_HS = "m_axi_rmem7_R.data" *)input m_axi_rmem7_RLAST;
  (* RS_HS = "m_axi_rmem7_R.ready" *)output m_axi_rmem7_RREADY;
  (* RS_HS = "m_axi_rmem7_R.data" *)input [1:0] m_axi_rmem7_RRESP;
  (* RS_HS = "m_axi_rmem7_R.valid" *)input m_axi_rmem7_RVALID;
  (* RS_HS = "m_axi_rmem7_W.data" *)output [511:0] m_axi_rmem7_WDATA;
  (* RS_HS = "m_axi_rmem7_W.data" *)output m_axi_rmem7_WLAST;
  (* RS_HS = "m_axi_rmem7_W.ready" *)input m_axi_rmem7_WREADY;
  (* RS_HS = "m_axi_rmem7_W.data" *)output [63:0] m_axi_rmem7_WSTRB;
  (* RS_HS = "m_axi_rmem7_W.valid" *)output m_axi_rmem7_WVALID;
  (* RS_HS = "m_axi_rmem8_AR.data" *)output [63:0] m_axi_rmem8_ARADDR;
  (* RS_HS = "m_axi_rmem8_AR.data" *)output [1:0] m_axi_rmem8_ARBURST;
  (* RS_HS = "m_axi_rmem8_AR.data" *)output [3:0] m_axi_rmem8_ARCACHE;
  (* RS_HS = "m_axi_rmem8_AR.data" *)output [1:0] m_axi_rmem8_ARID;
  (* RS_HS = "m_axi_rmem8_AR.data" *)output [7:0] m_axi_rmem8_ARLEN;
  (* RS_HS = "m_axi_rmem8_AR.data" *)output m_axi_rmem8_ARLOCK;
  (* RS_HS = "m_axi_rmem8_AR.data" *)output [2:0] m_axi_rmem8_ARPROT;
  (* RS_HS = "m_axi_rmem8_AR.data" *)output [3:0] m_axi_rmem8_ARQOS;
  (* RS_HS = "m_axi_rmem8_AR.ready" *)input m_axi_rmem8_ARREADY;
  (* RS_HS = "m_axi_rmem8_AR.data" *)output [2:0] m_axi_rmem8_ARSIZE;
  (* RS_HS = "m_axi_rmem8_AR.valid" *)output m_axi_rmem8_ARVALID;
  (* RS_HS = "m_axi_rmem8_AW.data" *)output [63:0] m_axi_rmem8_AWADDR;
  (* RS_HS = "m_axi_rmem8_AW.data" *)output [1:0] m_axi_rmem8_AWBURST;
  (* RS_HS = "m_axi_rmem8_AW.data" *)output [3:0] m_axi_rmem8_AWCACHE;
  (* RS_HS = "m_axi_rmem8_AW.data" *)output [1:0] m_axi_rmem8_AWID;
  (* RS_HS = "m_axi_rmem8_AW.data" *)output [7:0] m_axi_rmem8_AWLEN;
  (* RS_HS = "m_axi_rmem8_AW.data" *)output m_axi_rmem8_AWLOCK;
  (* RS_HS = "m_axi_rmem8_AW.data" *)output [2:0] m_axi_rmem8_AWPROT;
  (* RS_HS = "m_axi_rmem8_AW.data" *)output [3:0] m_axi_rmem8_AWQOS;
  (* RS_HS = "m_axi_rmem8_AW.ready" *)input m_axi_rmem8_AWREADY;
  (* RS_HS = "m_axi_rmem8_AW.data" *)output [2:0] m_axi_rmem8_AWSIZE;
  (* RS_HS = "m_axi_rmem8_AW.valid" *)output m_axi_rmem8_AWVALID;
  (* RS_HS = "m_axi_rmem8_B.data" *)input [1:0] m_axi_rmem8_BID;
  (* RS_HS = "m_axi_rmem8_B.ready" *)output m_axi_rmem8_BREADY;
  (* RS_HS = "m_axi_rmem8_B.data" *)input [1:0] m_axi_rmem8_BRESP;
  (* RS_HS = "m_axi_rmem8_B.valid" *)input m_axi_rmem8_BVALID;
  (* RS_HS = "m_axi_rmem8_R.data" *)input [511:0] m_axi_rmem8_RDATA;
  (* RS_HS = "m_axi_rmem8_R.data" *)input [1:0] m_axi_rmem8_RID;
  (* RS_HS = "m_axi_rmem8_R.data" *)input m_axi_rmem8_RLAST;
  (* RS_HS = "m_axi_rmem8_R.ready" *)output m_axi_rmem8_RREADY;
  (* RS_HS = "m_axi_rmem8_R.data" *)input [1:0] m_axi_rmem8_RRESP;
  (* RS_HS = "m_axi_rmem8_R.valid" *)input m_axi_rmem8_RVALID;
  (* RS_HS = "m_axi_rmem8_W.data" *)output [511:0] m_axi_rmem8_WDATA;
  (* RS_HS = "m_axi_rmem8_W.data" *)output m_axi_rmem8_WLAST;
  (* RS_HS = "m_axi_rmem8_W.ready" *)input m_axi_rmem8_WREADY;
  (* RS_HS = "m_axi_rmem8_W.data" *)output [63:0] m_axi_rmem8_WSTRB;
  (* RS_HS = "m_axi_rmem8_W.valid" *)output m_axi_rmem8_WVALID;
  (* RS_HS = "m_axi_rmem9_AR.data" *)output [63:0] m_axi_rmem9_ARADDR;
  (* RS_HS = "m_axi_rmem9_AR.data" *)output [1:0] m_axi_rmem9_ARBURST;
  (* RS_HS = "m_axi_rmem9_AR.data" *)output [3:0] m_axi_rmem9_ARCACHE;
  (* RS_HS = "m_axi_rmem9_AR.data" *)output [1:0] m_axi_rmem9_ARID;
  (* RS_HS = "m_axi_rmem9_AR.data" *)output [7:0] m_axi_rmem9_ARLEN;
  (* RS_HS = "m_axi_rmem9_AR.data" *)output m_axi_rmem9_ARLOCK;
  (* RS_HS = "m_axi_rmem9_AR.data" *)output [2:0] m_axi_rmem9_ARPROT;
  (* RS_HS = "m_axi_rmem9_AR.data" *)output [3:0] m_axi_rmem9_ARQOS;
  (* RS_HS = "m_axi_rmem9_AR.ready" *)input m_axi_rmem9_ARREADY;
  (* RS_HS = "m_axi_rmem9_AR.data" *)output [2:0] m_axi_rmem9_ARSIZE;
  (* RS_HS = "m_axi_rmem9_AR.valid" *)output m_axi_rmem9_ARVALID;
  (* RS_HS = "m_axi_rmem9_AW.data" *)output [63:0] m_axi_rmem9_AWADDR;
  (* RS_HS = "m_axi_rmem9_AW.data" *)output [1:0] m_axi_rmem9_AWBURST;
  (* RS_HS = "m_axi_rmem9_AW.data" *)output [3:0] m_axi_rmem9_AWCACHE;
  (* RS_HS = "m_axi_rmem9_AW.data" *)output [1:0] m_axi_rmem9_AWID;
  (* RS_HS = "m_axi_rmem9_AW.data" *)output [7:0] m_axi_rmem9_AWLEN;
  (* RS_HS = "m_axi_rmem9_AW.data" *)output m_axi_rmem9_AWLOCK;
  (* RS_HS = "m_axi_rmem9_AW.data" *)output [2:0] m_axi_rmem9_AWPROT;
  (* RS_HS = "m_axi_rmem9_AW.data" *)output [3:0] m_axi_rmem9_AWQOS;
  (* RS_HS = "m_axi_rmem9_AW.ready" *)input m_axi_rmem9_AWREADY;
  (* RS_HS = "m_axi_rmem9_AW.data" *)output [2:0] m_axi_rmem9_AWSIZE;
  (* RS_HS = "m_axi_rmem9_AW.valid" *)output m_axi_rmem9_AWVALID;
  (* RS_HS = "m_axi_rmem9_B.data" *)input [1:0] m_axi_rmem9_BID;
  (* RS_HS = "m_axi_rmem9_B.ready" *)output m_axi_rmem9_BREADY;
  (* RS_HS = "m_axi_rmem9_B.data" *)input [1:0] m_axi_rmem9_BRESP;
  (* RS_HS = "m_axi_rmem9_B.valid" *)input m_axi_rmem9_BVALID;
  (* RS_HS = "m_axi_rmem9_R.data" *)input [511:0] m_axi_rmem9_RDATA;
  (* RS_HS = "m_axi_rmem9_R.data" *)input [1:0] m_axi_rmem9_RID;
  (* RS_HS = "m_axi_rmem9_R.data" *)input m_axi_rmem9_RLAST;
  (* RS_HS = "m_axi_rmem9_R.ready" *)output m_axi_rmem9_RREADY;
  (* RS_HS = "m_axi_rmem9_R.data" *)input [1:0] m_axi_rmem9_RRESP;
  (* RS_HS = "m_axi_rmem9_R.valid" *)input m_axi_rmem9_RVALID;
  (* RS_HS = "m_axi_rmem9_W.data" *)output [511:0] m_axi_rmem9_WDATA;
  (* RS_HS = "m_axi_rmem9_W.data" *)output m_axi_rmem9_WLAST;
  (* RS_HS = "m_axi_rmem9_W.ready" *)input m_axi_rmem9_WREADY;
  (* RS_HS = "m_axi_rmem9_W.data" *)output [63:0] m_axi_rmem9_WSTRB;
  (* RS_HS = "m_axi_rmem9_W.valid" *)output m_axi_rmem9_WVALID;
  (* RS_HS = "m_axi_rmem10_AR.data" *)output [63:0] m_axi_rmem10_ARADDR;
  (* RS_HS = "m_axi_rmem10_AR.data" *)output [1:0] m_axi_rmem10_ARBURST;
  (* RS_HS = "m_axi_rmem10_AR.data" *)output [3:0] m_axi_rmem10_ARCACHE;
  (* RS_HS = "m_axi_rmem10_AR.data" *)output [1:0] m_axi_rmem10_ARID;
  (* RS_HS = "m_axi_rmem10_AR.data" *)output [7:0] m_axi_rmem10_ARLEN;
  (* RS_HS = "m_axi_rmem10_AR.data" *)output m_axi_rmem10_ARLOCK;
  (* RS_HS = "m_axi_rmem10_AR.data" *)output [2:0] m_axi_rmem10_ARPROT;
  (* RS_HS = "m_axi_rmem10_AR.data" *)output [3:0] m_axi_rmem10_ARQOS;
  (* RS_HS = "m_axi_rmem10_AR.ready" *)input m_axi_rmem10_ARREADY;
  (* RS_HS = "m_axi_rmem10_AR.data" *)output [2:0] m_axi_rmem10_ARSIZE;
  (* RS_HS = "m_axi_rmem10_AR.valid" *)output m_axi_rmem10_ARVALID;
  (* RS_HS = "m_axi_rmem10_AW.data" *)output [63:0] m_axi_rmem10_AWADDR;
  (* RS_HS = "m_axi_rmem10_AW.data" *)output [1:0] m_axi_rmem10_AWBURST;
  (* RS_HS = "m_axi_rmem10_AW.data" *)output [3:0] m_axi_rmem10_AWCACHE;
  (* RS_HS = "m_axi_rmem10_AW.data" *)output [1:0] m_axi_rmem10_AWID;
  (* RS_HS = "m_axi_rmem10_AW.data" *)output [7:0] m_axi_rmem10_AWLEN;
  (* RS_HS = "m_axi_rmem10_AW.data" *)output m_axi_rmem10_AWLOCK;
  (* RS_HS = "m_axi_rmem10_AW.data" *)output [2:0] m_axi_rmem10_AWPROT;
  (* RS_HS = "m_axi_rmem10_AW.data" *)output [3:0] m_axi_rmem10_AWQOS;
  (* RS_HS = "m_axi_rmem10_AW.ready" *)input m_axi_rmem10_AWREADY;
  (* RS_HS = "m_axi_rmem10_AW.data" *)output [2:0] m_axi_rmem10_AWSIZE;
  (* RS_HS = "m_axi_rmem10_AW.valid" *)output m_axi_rmem10_AWVALID;
  (* RS_HS = "m_axi_rmem10_B.data" *)input [1:0] m_axi_rmem10_BID;
  (* RS_HS = "m_axi_rmem10_B.ready" *)output m_axi_rmem10_BREADY;
  (* RS_HS = "m_axi_rmem10_B.data" *)input [1:0] m_axi_rmem10_BRESP;
  (* RS_HS = "m_axi_rmem10_B.valid" *)input m_axi_rmem10_BVALID;
  (* RS_HS = "m_axi_rmem10_R.data" *)input [511:0] m_axi_rmem10_RDATA;
  (* RS_HS = "m_axi_rmem10_R.data" *)input [1:0] m_axi_rmem10_RID;
  (* RS_HS = "m_axi_rmem10_R.data" *)input m_axi_rmem10_RLAST;
  (* RS_HS = "m_axi_rmem10_R.ready" *)output m_axi_rmem10_RREADY;
  (* RS_HS = "m_axi_rmem10_R.data" *)input [1:0] m_axi_rmem10_RRESP;
  (* RS_HS = "m_axi_rmem10_R.valid" *)input m_axi_rmem10_RVALID;
  (* RS_HS = "m_axi_rmem10_W.data" *)output [511:0] m_axi_rmem10_WDATA;
  (* RS_HS = "m_axi_rmem10_W.data" *)output m_axi_rmem10_WLAST;
  (* RS_HS = "m_axi_rmem10_W.ready" *)input m_axi_rmem10_WREADY;
  (* RS_HS = "m_axi_rmem10_W.data" *)output [63:0] m_axi_rmem10_WSTRB;
  (* RS_HS = "m_axi_rmem10_W.valid" *)output m_axi_rmem10_WVALID;
  (* RS_HS = "m_axi_rmem11_AR.data" *)output [63:0] m_axi_rmem11_ARADDR;
  (* RS_HS = "m_axi_rmem11_AR.data" *)output [1:0] m_axi_rmem11_ARBURST;
  (* RS_HS = "m_axi_rmem11_AR.data" *)output [3:0] m_axi_rmem11_ARCACHE;
  (* RS_HS = "m_axi_rmem11_AR.data" *)output [1:0] m_axi_rmem11_ARID;
  (* RS_HS = "m_axi_rmem11_AR.data" *)output [7:0] m_axi_rmem11_ARLEN;
  (* RS_HS = "m_axi_rmem11_AR.data" *)output m_axi_rmem11_ARLOCK;
  (* RS_HS = "m_axi_rmem11_AR.data" *)output [2:0] m_axi_rmem11_ARPROT;
  (* RS_HS = "m_axi_rmem11_AR.data" *)output [3:0] m_axi_rmem11_ARQOS;
  (* RS_HS = "m_axi_rmem11_AR.ready" *)input m_axi_rmem11_ARREADY;
  (* RS_HS = "m_axi_rmem11_AR.data" *)output [2:0] m_axi_rmem11_ARSIZE;
  (* RS_HS = "m_axi_rmem11_AR.valid" *)output m_axi_rmem11_ARVALID;
  (* RS_HS = "m_axi_rmem11_AW.data" *)output [63:0] m_axi_rmem11_AWADDR;
  (* RS_HS = "m_axi_rmem11_AW.data" *)output [1:0] m_axi_rmem11_AWBURST;
  (* RS_HS = "m_axi_rmem11_AW.data" *)output [3:0] m_axi_rmem11_AWCACHE;
  (* RS_HS = "m_axi_rmem11_AW.data" *)output [1:0] m_axi_rmem11_AWID;
  (* RS_HS = "m_axi_rmem11_AW.data" *)output [7:0] m_axi_rmem11_AWLEN;
  (* RS_HS = "m_axi_rmem11_AW.data" *)output m_axi_rmem11_AWLOCK;
  (* RS_HS = "m_axi_rmem11_AW.data" *)output [2:0] m_axi_rmem11_AWPROT;
  (* RS_HS = "m_axi_rmem11_AW.data" *)output [3:0] m_axi_rmem11_AWQOS;
  (* RS_HS = "m_axi_rmem11_AW.ready" *)input m_axi_rmem11_AWREADY;
  (* RS_HS = "m_axi_rmem11_AW.data" *)output [2:0] m_axi_rmem11_AWSIZE;
  (* RS_HS = "m_axi_rmem11_AW.valid" *)output m_axi_rmem11_AWVALID;
  (* RS_HS = "m_axi_rmem11_B.data" *)input [1:0] m_axi_rmem11_BID;
  (* RS_HS = "m_axi_rmem11_B.ready" *)output m_axi_rmem11_BREADY;
  (* RS_HS = "m_axi_rmem11_B.data" *)input [1:0] m_axi_rmem11_BRESP;
  (* RS_HS = "m_axi_rmem11_B.valid" *)input m_axi_rmem11_BVALID;
  (* RS_HS = "m_axi_rmem11_R.data" *)input [511:0] m_axi_rmem11_RDATA;
  (* RS_HS = "m_axi_rmem11_R.data" *)input [1:0] m_axi_rmem11_RID;
  (* RS_HS = "m_axi_rmem11_R.data" *)input m_axi_rmem11_RLAST;
  (* RS_HS = "m_axi_rmem11_R.ready" *)output m_axi_rmem11_RREADY;
  (* RS_HS = "m_axi_rmem11_R.data" *)input [1:0] m_axi_rmem11_RRESP;
  (* RS_HS = "m_axi_rmem11_R.valid" *)input m_axi_rmem11_RVALID;
  (* RS_HS = "m_axi_rmem11_W.data" *)output [511:0] m_axi_rmem11_WDATA;
  (* RS_HS = "m_axi_rmem11_W.data" *)output m_axi_rmem11_WLAST;
  (* RS_HS = "m_axi_rmem11_W.ready" *)input m_axi_rmem11_WREADY;
  (* RS_HS = "m_axi_rmem11_W.data" *)output [63:0] m_axi_rmem11_WSTRB;
  (* RS_HS = "m_axi_rmem11_W.valid" *)output m_axi_rmem11_WVALID;
  (* RS_HS = "m_axi_rmem12_AR.data" *)output [63:0] m_axi_rmem12_ARADDR;
  (* RS_HS = "m_axi_rmem12_AR.data" *)output [1:0] m_axi_rmem12_ARBURST;
  (* RS_HS = "m_axi_rmem12_AR.data" *)output [3:0] m_axi_rmem12_ARCACHE;
  (* RS_HS = "m_axi_rmem12_AR.data" *)output [1:0] m_axi_rmem12_ARID;
  (* RS_HS = "m_axi_rmem12_AR.data" *)output [7:0] m_axi_rmem12_ARLEN;
  (* RS_HS = "m_axi_rmem12_AR.data" *)output m_axi_rmem12_ARLOCK;
  (* RS_HS = "m_axi_rmem12_AR.data" *)output [2:0] m_axi_rmem12_ARPROT;
  (* RS_HS = "m_axi_rmem12_AR.data" *)output [3:0] m_axi_rmem12_ARQOS;
  (* RS_HS = "m_axi_rmem12_AR.ready" *)input m_axi_rmem12_ARREADY;
  (* RS_HS = "m_axi_rmem12_AR.data" *)output [2:0] m_axi_rmem12_ARSIZE;
  (* RS_HS = "m_axi_rmem12_AR.valid" *)output m_axi_rmem12_ARVALID;
  (* RS_HS = "m_axi_rmem12_AW.data" *)output [63:0] m_axi_rmem12_AWADDR;
  (* RS_HS = "m_axi_rmem12_AW.data" *)output [1:0] m_axi_rmem12_AWBURST;
  (* RS_HS = "m_axi_rmem12_AW.data" *)output [3:0] m_axi_rmem12_AWCACHE;
  (* RS_HS = "m_axi_rmem12_AW.data" *)output [1:0] m_axi_rmem12_AWID;
  (* RS_HS = "m_axi_rmem12_AW.data" *)output [7:0] m_axi_rmem12_AWLEN;
  (* RS_HS = "m_axi_rmem12_AW.data" *)output m_axi_rmem12_AWLOCK;
  (* RS_HS = "m_axi_rmem12_AW.data" *)output [2:0] m_axi_rmem12_AWPROT;
  (* RS_HS = "m_axi_rmem12_AW.data" *)output [3:0] m_axi_rmem12_AWQOS;
  (* RS_HS = "m_axi_rmem12_AW.ready" *)input m_axi_rmem12_AWREADY;
  (* RS_HS = "m_axi_rmem12_AW.data" *)output [2:0] m_axi_rmem12_AWSIZE;
  (* RS_HS = "m_axi_rmem12_AW.valid" *)output m_axi_rmem12_AWVALID;
  (* RS_HS = "m_axi_rmem12_B.data" *)input [1:0] m_axi_rmem12_BID;
  (* RS_HS = "m_axi_rmem12_B.ready" *)output m_axi_rmem12_BREADY;
  (* RS_HS = "m_axi_rmem12_B.data" *)input [1:0] m_axi_rmem12_BRESP;
  (* RS_HS = "m_axi_rmem12_B.valid" *)input m_axi_rmem12_BVALID;
  (* RS_HS = "m_axi_rmem12_R.data" *)input [511:0] m_axi_rmem12_RDATA;
  (* RS_HS = "m_axi_rmem12_R.data" *)input [1:0] m_axi_rmem12_RID;
  (* RS_HS = "m_axi_rmem12_R.data" *)input m_axi_rmem12_RLAST;
  (* RS_HS = "m_axi_rmem12_R.ready" *)output m_axi_rmem12_RREADY;
  (* RS_HS = "m_axi_rmem12_R.data" *)input [1:0] m_axi_rmem12_RRESP;
  (* RS_HS = "m_axi_rmem12_R.valid" *)input m_axi_rmem12_RVALID;
  (* RS_HS = "m_axi_rmem12_W.data" *)output [511:0] m_axi_rmem12_WDATA;
  (* RS_HS = "m_axi_rmem12_W.data" *)output m_axi_rmem12_WLAST;
  (* RS_HS = "m_axi_rmem12_W.ready" *)input m_axi_rmem12_WREADY;
  (* RS_HS = "m_axi_rmem12_W.data" *)output [63:0] m_axi_rmem12_WSTRB;
  (* RS_HS = "m_axi_rmem12_W.valid" *)output m_axi_rmem12_WVALID;
  (* RS_HS = "m_axi_rmem13_AR.data" *)output [63:0] m_axi_rmem13_ARADDR;
  (* RS_HS = "m_axi_rmem13_AR.data" *)output [1:0] m_axi_rmem13_ARBURST;
  (* RS_HS = "m_axi_rmem13_AR.data" *)output [3:0] m_axi_rmem13_ARCACHE;
  (* RS_HS = "m_axi_rmem13_AR.data" *)output [1:0] m_axi_rmem13_ARID;
  (* RS_HS = "m_axi_rmem13_AR.data" *)output [7:0] m_axi_rmem13_ARLEN;
  (* RS_HS = "m_axi_rmem13_AR.data" *)output m_axi_rmem13_ARLOCK;
  (* RS_HS = "m_axi_rmem13_AR.data" *)output [2:0] m_axi_rmem13_ARPROT;
  (* RS_HS = "m_axi_rmem13_AR.data" *)output [3:0] m_axi_rmem13_ARQOS;
  (* RS_HS = "m_axi_rmem13_AR.ready" *)input m_axi_rmem13_ARREADY;
  (* RS_HS = "m_axi_rmem13_AR.data" *)output [2:0] m_axi_rmem13_ARSIZE;
  (* RS_HS = "m_axi_rmem13_AR.valid" *)output m_axi_rmem13_ARVALID;
  (* RS_HS = "m_axi_rmem13_AW.data" *)output [63:0] m_axi_rmem13_AWADDR;
  (* RS_HS = "m_axi_rmem13_AW.data" *)output [1:0] m_axi_rmem13_AWBURST;
  (* RS_HS = "m_axi_rmem13_AW.data" *)output [3:0] m_axi_rmem13_AWCACHE;
  (* RS_HS = "m_axi_rmem13_AW.data" *)output [1:0] m_axi_rmem13_AWID;
  (* RS_HS = "m_axi_rmem13_AW.data" *)output [7:0] m_axi_rmem13_AWLEN;
  (* RS_HS = "m_axi_rmem13_AW.data" *)output m_axi_rmem13_AWLOCK;
  (* RS_HS = "m_axi_rmem13_AW.data" *)output [2:0] m_axi_rmem13_AWPROT;
  (* RS_HS = "m_axi_rmem13_AW.data" *)output [3:0] m_axi_rmem13_AWQOS;
  (* RS_HS = "m_axi_rmem13_AW.ready" *)input m_axi_rmem13_AWREADY;
  (* RS_HS = "m_axi_rmem13_AW.data" *)output [2:0] m_axi_rmem13_AWSIZE;
  (* RS_HS = "m_axi_rmem13_AW.valid" *)output m_axi_rmem13_AWVALID;
  (* RS_HS = "m_axi_rmem13_B.data" *)input [1:0] m_axi_rmem13_BID;
  (* RS_HS = "m_axi_rmem13_B.ready" *)output m_axi_rmem13_BREADY;
  (* RS_HS = "m_axi_rmem13_B.data" *)input [1:0] m_axi_rmem13_BRESP;
  (* RS_HS = "m_axi_rmem13_B.valid" *)input m_axi_rmem13_BVALID;
  (* RS_HS = "m_axi_rmem13_R.data" *)input [511:0] m_axi_rmem13_RDATA;
  (* RS_HS = "m_axi_rmem13_R.data" *)input [1:0] m_axi_rmem13_RID;
  (* RS_HS = "m_axi_rmem13_R.data" *)input m_axi_rmem13_RLAST;
  (* RS_HS = "m_axi_rmem13_R.ready" *)output m_axi_rmem13_RREADY;
  (* RS_HS = "m_axi_rmem13_R.data" *)input [1:0] m_axi_rmem13_RRESP;
  (* RS_HS = "m_axi_rmem13_R.valid" *)input m_axi_rmem13_RVALID;
  (* RS_HS = "m_axi_rmem13_W.data" *)output [511:0] m_axi_rmem13_WDATA;
  (* RS_HS = "m_axi_rmem13_W.data" *)output m_axi_rmem13_WLAST;
  (* RS_HS = "m_axi_rmem13_W.ready" *)input m_axi_rmem13_WREADY;
  (* RS_HS = "m_axi_rmem13_W.data" *)output [63:0] m_axi_rmem13_WSTRB;
  (* RS_HS = "m_axi_rmem13_W.valid" *)output m_axi_rmem13_WVALID;
  (* RS_HS = "m_axi_rmem14_AR.data" *)output [63:0] m_axi_rmem14_ARADDR;
  (* RS_HS = "m_axi_rmem14_AR.data" *)output [1:0] m_axi_rmem14_ARBURST;
  (* RS_HS = "m_axi_rmem14_AR.data" *)output [3:0] m_axi_rmem14_ARCACHE;
  (* RS_HS = "m_axi_rmem14_AR.data" *)output [1:0] m_axi_rmem14_ARID;
  (* RS_HS = "m_axi_rmem14_AR.data" *)output [7:0] m_axi_rmem14_ARLEN;
  (* RS_HS = "m_axi_rmem14_AR.data" *)output m_axi_rmem14_ARLOCK;
  (* RS_HS = "m_axi_rmem14_AR.data" *)output [2:0] m_axi_rmem14_ARPROT;
  (* RS_HS = "m_axi_rmem14_AR.data" *)output [3:0] m_axi_rmem14_ARQOS;
  (* RS_HS = "m_axi_rmem14_AR.ready" *)input m_axi_rmem14_ARREADY;
  (* RS_HS = "m_axi_rmem14_AR.data" *)output [2:0] m_axi_rmem14_ARSIZE;
  (* RS_HS = "m_axi_rmem14_AR.valid" *)output m_axi_rmem14_ARVALID;
  (* RS_HS = "m_axi_rmem14_AW.data" *)output [63:0] m_axi_rmem14_AWADDR;
  (* RS_HS = "m_axi_rmem14_AW.data" *)output [1:0] m_axi_rmem14_AWBURST;
  (* RS_HS = "m_axi_rmem14_AW.data" *)output [3:0] m_axi_rmem14_AWCACHE;
  (* RS_HS = "m_axi_rmem14_AW.data" *)output [1:0] m_axi_rmem14_AWID;
  (* RS_HS = "m_axi_rmem14_AW.data" *)output [7:0] m_axi_rmem14_AWLEN;
  (* RS_HS = "m_axi_rmem14_AW.data" *)output m_axi_rmem14_AWLOCK;
  (* RS_HS = "m_axi_rmem14_AW.data" *)output [2:0] m_axi_rmem14_AWPROT;
  (* RS_HS = "m_axi_rmem14_AW.data" *)output [3:0] m_axi_rmem14_AWQOS;
  (* RS_HS = "m_axi_rmem14_AW.ready" *)input m_axi_rmem14_AWREADY;
  (* RS_HS = "m_axi_rmem14_AW.data" *)output [2:0] m_axi_rmem14_AWSIZE;
  (* RS_HS = "m_axi_rmem14_AW.valid" *)output m_axi_rmem14_AWVALID;
  (* RS_HS = "m_axi_rmem14_B.data" *)input [1:0] m_axi_rmem14_BID;
  (* RS_HS = "m_axi_rmem14_B.ready" *)output m_axi_rmem14_BREADY;
  (* RS_HS = "m_axi_rmem14_B.data" *)input [1:0] m_axi_rmem14_BRESP;
  (* RS_HS = "m_axi_rmem14_B.valid" *)input m_axi_rmem14_BVALID;
  (* RS_HS = "m_axi_rmem14_R.data" *)input [511:0] m_axi_rmem14_RDATA;
  (* RS_HS = "m_axi_rmem14_R.data" *)input [1:0] m_axi_rmem14_RID;
  (* RS_HS = "m_axi_rmem14_R.data" *)input m_axi_rmem14_RLAST;
  (* RS_HS = "m_axi_rmem14_R.ready" *)output m_axi_rmem14_RREADY;
  (* RS_HS = "m_axi_rmem14_R.data" *)input [1:0] m_axi_rmem14_RRESP;
  (* RS_HS = "m_axi_rmem14_R.valid" *)input m_axi_rmem14_RVALID;
  (* RS_HS = "m_axi_rmem14_W.data" *)output [511:0] m_axi_rmem14_WDATA;
  (* RS_HS = "m_axi_rmem14_W.data" *)output m_axi_rmem14_WLAST;
  (* RS_HS = "m_axi_rmem14_W.ready" *)input m_axi_rmem14_WREADY;
  (* RS_HS = "m_axi_rmem14_W.data" *)output [63:0] m_axi_rmem14_WSTRB;
  (* RS_HS = "m_axi_rmem14_W.valid" *)output m_axi_rmem14_WVALID;
  (* RS_HS = "m_axi_rmem15_AR.data" *)output [63:0] m_axi_rmem15_ARADDR;
  (* RS_HS = "m_axi_rmem15_AR.data" *)output [1:0] m_axi_rmem15_ARBURST;
  (* RS_HS = "m_axi_rmem15_AR.data" *)output [3:0] m_axi_rmem15_ARCACHE;
  (* RS_HS = "m_axi_rmem15_AR.data" *)output [1:0] m_axi_rmem15_ARID;
  (* RS_HS = "m_axi_rmem15_AR.data" *)output [7:0] m_axi_rmem15_ARLEN;
  (* RS_HS = "m_axi_rmem15_AR.data" *)output m_axi_rmem15_ARLOCK;
  (* RS_HS = "m_axi_rmem15_AR.data" *)output [2:0] m_axi_rmem15_ARPROT;
  (* RS_HS = "m_axi_rmem15_AR.data" *)output [3:0] m_axi_rmem15_ARQOS;
  (* RS_HS = "m_axi_rmem15_AR.ready" *)input m_axi_rmem15_ARREADY;
  (* RS_HS = "m_axi_rmem15_AR.data" *)output [2:0] m_axi_rmem15_ARSIZE;
  (* RS_HS = "m_axi_rmem15_AR.valid" *)output m_axi_rmem15_ARVALID;
  (* RS_HS = "m_axi_rmem15_AW.data" *)output [63:0] m_axi_rmem15_AWADDR;
  (* RS_HS = "m_axi_rmem15_AW.data" *)output [1:0] m_axi_rmem15_AWBURST;
  (* RS_HS = "m_axi_rmem15_AW.data" *)output [3:0] m_axi_rmem15_AWCACHE;
  (* RS_HS = "m_axi_rmem15_AW.data" *)output [1:0] m_axi_rmem15_AWID;
  (* RS_HS = "m_axi_rmem15_AW.data" *)output [7:0] m_axi_rmem15_AWLEN;
  (* RS_HS = "m_axi_rmem15_AW.data" *)output m_axi_rmem15_AWLOCK;
  (* RS_HS = "m_axi_rmem15_AW.data" *)output [2:0] m_axi_rmem15_AWPROT;
  (* RS_HS = "m_axi_rmem15_AW.data" *)output [3:0] m_axi_rmem15_AWQOS;
  (* RS_HS = "m_axi_rmem15_AW.ready" *)input m_axi_rmem15_AWREADY;
  (* RS_HS = "m_axi_rmem15_AW.data" *)output [2:0] m_axi_rmem15_AWSIZE;
  (* RS_HS = "m_axi_rmem15_AW.valid" *)output m_axi_rmem15_AWVALID;
  (* RS_HS = "m_axi_rmem15_B.data" *)input [1:0] m_axi_rmem15_BID;
  (* RS_HS = "m_axi_rmem15_B.ready" *)output m_axi_rmem15_BREADY;
  (* RS_HS = "m_axi_rmem15_B.data" *)input [1:0] m_axi_rmem15_BRESP;
  (* RS_HS = "m_axi_rmem15_B.valid" *)input m_axi_rmem15_BVALID;
  (* RS_HS = "m_axi_rmem15_R.data" *)input [511:0] m_axi_rmem15_RDATA;
  (* RS_HS = "m_axi_rmem15_R.data" *)input [1:0] m_axi_rmem15_RID;
  (* RS_HS = "m_axi_rmem15_R.data" *)input m_axi_rmem15_RLAST;
  (* RS_HS = "m_axi_rmem15_R.ready" *)output m_axi_rmem15_RREADY;
  (* RS_HS = "m_axi_rmem15_R.data" *)input [1:0] m_axi_rmem15_RRESP;
  (* RS_HS = "m_axi_rmem15_R.valid" *)input m_axi_rmem15_RVALID;
  (* RS_HS = "m_axi_rmem15_W.data" *)output [511:0] m_axi_rmem15_WDATA;
  (* RS_HS = "m_axi_rmem15_W.data" *)output m_axi_rmem15_WLAST;
  (* RS_HS = "m_axi_rmem15_W.ready" *)input m_axi_rmem15_WREADY;
  (* RS_HS = "m_axi_rmem15_W.data" *)output [63:0] m_axi_rmem15_WSTRB;
  (* RS_HS = "m_axi_rmem15_W.valid" *)output m_axi_rmem15_WVALID;
  (* RS_HS = "m_axi_rmem16_AR.data" *)output [63:0] m_axi_rmem16_ARADDR;
  (* RS_HS = "m_axi_rmem16_AR.data" *)output [1:0] m_axi_rmem16_ARBURST;
  (* RS_HS = "m_axi_rmem16_AR.data" *)output [3:0] m_axi_rmem16_ARCACHE;
  (* RS_HS = "m_axi_rmem16_AR.data" *)output [1:0] m_axi_rmem16_ARID;
  (* RS_HS = "m_axi_rmem16_AR.data" *)output [7:0] m_axi_rmem16_ARLEN;
  (* RS_HS = "m_axi_rmem16_AR.data" *)output m_axi_rmem16_ARLOCK;
  (* RS_HS = "m_axi_rmem16_AR.data" *)output [2:0] m_axi_rmem16_ARPROT;
  (* RS_HS = "m_axi_rmem16_AR.data" *)output [3:0] m_axi_rmem16_ARQOS;
  (* RS_HS = "m_axi_rmem16_AR.ready" *)input m_axi_rmem16_ARREADY;
  (* RS_HS = "m_axi_rmem16_AR.data" *)output [2:0] m_axi_rmem16_ARSIZE;
  (* RS_HS = "m_axi_rmem16_AR.valid" *)output m_axi_rmem16_ARVALID;
  (* RS_HS = "m_axi_rmem16_AW.data" *)output [63:0] m_axi_rmem16_AWADDR;
  (* RS_HS = "m_axi_rmem16_AW.data" *)output [1:0] m_axi_rmem16_AWBURST;
  (* RS_HS = "m_axi_rmem16_AW.data" *)output [3:0] m_axi_rmem16_AWCACHE;
  (* RS_HS = "m_axi_rmem16_AW.data" *)output [1:0] m_axi_rmem16_AWID;
  (* RS_HS = "m_axi_rmem16_AW.data" *)output [7:0] m_axi_rmem16_AWLEN;
  (* RS_HS = "m_axi_rmem16_AW.data" *)output m_axi_rmem16_AWLOCK;
  (* RS_HS = "m_axi_rmem16_AW.data" *)output [2:0] m_axi_rmem16_AWPROT;
  (* RS_HS = "m_axi_rmem16_AW.data" *)output [3:0] m_axi_rmem16_AWQOS;
  (* RS_HS = "m_axi_rmem16_AW.ready" *)input m_axi_rmem16_AWREADY;
  (* RS_HS = "m_axi_rmem16_AW.data" *)output [2:0] m_axi_rmem16_AWSIZE;
  (* RS_HS = "m_axi_rmem16_AW.valid" *)output m_axi_rmem16_AWVALID;
  (* RS_HS = "m_axi_rmem16_B.data" *)input [1:0] m_axi_rmem16_BID;
  (* RS_HS = "m_axi_rmem16_B.ready" *)output m_axi_rmem16_BREADY;
  (* RS_HS = "m_axi_rmem16_B.data" *)input [1:0] m_axi_rmem16_BRESP;
  (* RS_HS = "m_axi_rmem16_B.valid" *)input m_axi_rmem16_BVALID;
  (* RS_HS = "m_axi_rmem16_R.data" *)input [511:0] m_axi_rmem16_RDATA;
  (* RS_HS = "m_axi_rmem16_R.data" *)input [1:0] m_axi_rmem16_RID;
  (* RS_HS = "m_axi_rmem16_R.data" *)input m_axi_rmem16_RLAST;
  (* RS_HS = "m_axi_rmem16_R.ready" *)output m_axi_rmem16_RREADY;
  (* RS_HS = "m_axi_rmem16_R.data" *)input [1:0] m_axi_rmem16_RRESP;
  (* RS_HS = "m_axi_rmem16_R.valid" *)input m_axi_rmem16_RVALID;
  (* RS_HS = "m_axi_rmem16_W.data" *)output [511:0] m_axi_rmem16_WDATA;
  (* RS_HS = "m_axi_rmem16_W.data" *)output m_axi_rmem16_WLAST;
  (* RS_HS = "m_axi_rmem16_W.ready" *)input m_axi_rmem16_WREADY;
  (* RS_HS = "m_axi_rmem16_W.data" *)output [63:0] m_axi_rmem16_WSTRB;
  (* RS_HS = "m_axi_rmem16_W.valid" *)output m_axi_rmem16_WVALID;
  (* RS_HS = "m_axi_rmem17_AR.data" *)output [63:0] m_axi_rmem17_ARADDR;
  (* RS_HS = "m_axi_rmem17_AR.data" *)output [1:0] m_axi_rmem17_ARBURST;
  (* RS_HS = "m_axi_rmem17_AR.data" *)output [3:0] m_axi_rmem17_ARCACHE;
  (* RS_HS = "m_axi_rmem17_AR.data" *)output [1:0] m_axi_rmem17_ARID;
  (* RS_HS = "m_axi_rmem17_AR.data" *)output [7:0] m_axi_rmem17_ARLEN;
  (* RS_HS = "m_axi_rmem17_AR.data" *)output m_axi_rmem17_ARLOCK;
  (* RS_HS = "m_axi_rmem17_AR.data" *)output [2:0] m_axi_rmem17_ARPROT;
  (* RS_HS = "m_axi_rmem17_AR.data" *)output [3:0] m_axi_rmem17_ARQOS;
  (* RS_HS = "m_axi_rmem17_AR.ready" *)input m_axi_rmem17_ARREADY;
  (* RS_HS = "m_axi_rmem17_AR.data" *)output [2:0] m_axi_rmem17_ARSIZE;
  (* RS_HS = "m_axi_rmem17_AR.valid" *)output m_axi_rmem17_ARVALID;
  (* RS_HS = "m_axi_rmem17_AW.data" *)output [63:0] m_axi_rmem17_AWADDR;
  (* RS_HS = "m_axi_rmem17_AW.data" *)output [1:0] m_axi_rmem17_AWBURST;
  (* RS_HS = "m_axi_rmem17_AW.data" *)output [3:0] m_axi_rmem17_AWCACHE;
  (* RS_HS = "m_axi_rmem17_AW.data" *)output [1:0] m_axi_rmem17_AWID;
  (* RS_HS = "m_axi_rmem17_AW.data" *)output [7:0] m_axi_rmem17_AWLEN;
  (* RS_HS = "m_axi_rmem17_AW.data" *)output m_axi_rmem17_AWLOCK;
  (* RS_HS = "m_axi_rmem17_AW.data" *)output [2:0] m_axi_rmem17_AWPROT;
  (* RS_HS = "m_axi_rmem17_AW.data" *)output [3:0] m_axi_rmem17_AWQOS;
  (* RS_HS = "m_axi_rmem17_AW.ready" *)input m_axi_rmem17_AWREADY;
  (* RS_HS = "m_axi_rmem17_AW.data" *)output [2:0] m_axi_rmem17_AWSIZE;
  (* RS_HS = "m_axi_rmem17_AW.valid" *)output m_axi_rmem17_AWVALID;
  (* RS_HS = "m_axi_rmem17_B.data" *)input [1:0] m_axi_rmem17_BID;
  (* RS_HS = "m_axi_rmem17_B.ready" *)output m_axi_rmem17_BREADY;
  (* RS_HS = "m_axi_rmem17_B.data" *)input [1:0] m_axi_rmem17_BRESP;
  (* RS_HS = "m_axi_rmem17_B.valid" *)input m_axi_rmem17_BVALID;
  (* RS_HS = "m_axi_rmem17_R.data" *)input [511:0] m_axi_rmem17_RDATA;
  (* RS_HS = "m_axi_rmem17_R.data" *)input [1:0] m_axi_rmem17_RID;
  (* RS_HS = "m_axi_rmem17_R.data" *)input m_axi_rmem17_RLAST;
  (* RS_HS = "m_axi_rmem17_R.ready" *)output m_axi_rmem17_RREADY;
  (* RS_HS = "m_axi_rmem17_R.data" *)input [1:0] m_axi_rmem17_RRESP;
  (* RS_HS = "m_axi_rmem17_R.valid" *)input m_axi_rmem17_RVALID;
  (* RS_HS = "m_axi_rmem17_W.data" *)output [511:0] m_axi_rmem17_WDATA;
  (* RS_HS = "m_axi_rmem17_W.data" *)output m_axi_rmem17_WLAST;
  (* RS_HS = "m_axi_rmem17_W.ready" *)input m_axi_rmem17_WREADY;
  (* RS_HS = "m_axi_rmem17_W.data" *)output [63:0] m_axi_rmem17_WSTRB;
  (* RS_HS = "m_axi_rmem17_W.valid" *)output m_axi_rmem17_WVALID;
  (* RS_HS = "m_axi_rmem18_AR.data" *)output [63:0] m_axi_rmem18_ARADDR;
  (* RS_HS = "m_axi_rmem18_AR.data" *)output [1:0] m_axi_rmem18_ARBURST;
  (* RS_HS = "m_axi_rmem18_AR.data" *)output [3:0] m_axi_rmem18_ARCACHE;
  (* RS_HS = "m_axi_rmem18_AR.data" *)output [1:0] m_axi_rmem18_ARID;
  (* RS_HS = "m_axi_rmem18_AR.data" *)output [7:0] m_axi_rmem18_ARLEN;
  (* RS_HS = "m_axi_rmem18_AR.data" *)output m_axi_rmem18_ARLOCK;
  (* RS_HS = "m_axi_rmem18_AR.data" *)output [2:0] m_axi_rmem18_ARPROT;
  (* RS_HS = "m_axi_rmem18_AR.data" *)output [3:0] m_axi_rmem18_ARQOS;
  (* RS_HS = "m_axi_rmem18_AR.ready" *)input m_axi_rmem18_ARREADY;
  (* RS_HS = "m_axi_rmem18_AR.data" *)output [2:0] m_axi_rmem18_ARSIZE;
  (* RS_HS = "m_axi_rmem18_AR.valid" *)output m_axi_rmem18_ARVALID;
  (* RS_HS = "m_axi_rmem18_AW.data" *)output [63:0] m_axi_rmem18_AWADDR;
  (* RS_HS = "m_axi_rmem18_AW.data" *)output [1:0] m_axi_rmem18_AWBURST;
  (* RS_HS = "m_axi_rmem18_AW.data" *)output [3:0] m_axi_rmem18_AWCACHE;
  (* RS_HS = "m_axi_rmem18_AW.data" *)output [1:0] m_axi_rmem18_AWID;
  (* RS_HS = "m_axi_rmem18_AW.data" *)output [7:0] m_axi_rmem18_AWLEN;
  (* RS_HS = "m_axi_rmem18_AW.data" *)output m_axi_rmem18_AWLOCK;
  (* RS_HS = "m_axi_rmem18_AW.data" *)output [2:0] m_axi_rmem18_AWPROT;
  (* RS_HS = "m_axi_rmem18_AW.data" *)output [3:0] m_axi_rmem18_AWQOS;
  (* RS_HS = "m_axi_rmem18_AW.ready" *)input m_axi_rmem18_AWREADY;
  (* RS_HS = "m_axi_rmem18_AW.data" *)output [2:0] m_axi_rmem18_AWSIZE;
  (* RS_HS = "m_axi_rmem18_AW.valid" *)output m_axi_rmem18_AWVALID;
  (* RS_HS = "m_axi_rmem18_B.data" *)input [1:0] m_axi_rmem18_BID;
  (* RS_HS = "m_axi_rmem18_B.ready" *)output m_axi_rmem18_BREADY;
  (* RS_HS = "m_axi_rmem18_B.data" *)input [1:0] m_axi_rmem18_BRESP;
  (* RS_HS = "m_axi_rmem18_B.valid" *)input m_axi_rmem18_BVALID;
  (* RS_HS = "m_axi_rmem18_R.data" *)input [511:0] m_axi_rmem18_RDATA;
  (* RS_HS = "m_axi_rmem18_R.data" *)input [1:0] m_axi_rmem18_RID;
  (* RS_HS = "m_axi_rmem18_R.data" *)input m_axi_rmem18_RLAST;
  (* RS_HS = "m_axi_rmem18_R.ready" *)output m_axi_rmem18_RREADY;
  (* RS_HS = "m_axi_rmem18_R.data" *)input [1:0] m_axi_rmem18_RRESP;
  (* RS_HS = "m_axi_rmem18_R.valid" *)input m_axi_rmem18_RVALID;
  (* RS_HS = "m_axi_rmem18_W.data" *)output [511:0] m_axi_rmem18_WDATA;
  (* RS_HS = "m_axi_rmem18_W.data" *)output m_axi_rmem18_WLAST;
  (* RS_HS = "m_axi_rmem18_W.ready" *)input m_axi_rmem18_WREADY;
  (* RS_HS = "m_axi_rmem18_W.data" *)output [63:0] m_axi_rmem18_WSTRB;
  (* RS_HS = "m_axi_rmem18_W.valid" *)output m_axi_rmem18_WVALID;
  (* RS_HS = "m_axi_rmem19_AR.data" *)output [63:0] m_axi_rmem19_ARADDR;
  (* RS_HS = "m_axi_rmem19_AR.data" *)output [1:0] m_axi_rmem19_ARBURST;
  (* RS_HS = "m_axi_rmem19_AR.data" *)output [3:0] m_axi_rmem19_ARCACHE;
  (* RS_HS = "m_axi_rmem19_AR.data" *)output [1:0] m_axi_rmem19_ARID;
  (* RS_HS = "m_axi_rmem19_AR.data" *)output [7:0] m_axi_rmem19_ARLEN;
  (* RS_HS = "m_axi_rmem19_AR.data" *)output m_axi_rmem19_ARLOCK;
  (* RS_HS = "m_axi_rmem19_AR.data" *)output [2:0] m_axi_rmem19_ARPROT;
  (* RS_HS = "m_axi_rmem19_AR.data" *)output [3:0] m_axi_rmem19_ARQOS;
  (* RS_HS = "m_axi_rmem19_AR.ready" *)input m_axi_rmem19_ARREADY;
  (* RS_HS = "m_axi_rmem19_AR.data" *)output [2:0] m_axi_rmem19_ARSIZE;
  (* RS_HS = "m_axi_rmem19_AR.valid" *)output m_axi_rmem19_ARVALID;
  (* RS_HS = "m_axi_rmem19_AW.data" *)output [63:0] m_axi_rmem19_AWADDR;
  (* RS_HS = "m_axi_rmem19_AW.data" *)output [1:0] m_axi_rmem19_AWBURST;
  (* RS_HS = "m_axi_rmem19_AW.data" *)output [3:0] m_axi_rmem19_AWCACHE;
  (* RS_HS = "m_axi_rmem19_AW.data" *)output [1:0] m_axi_rmem19_AWID;
  (* RS_HS = "m_axi_rmem19_AW.data" *)output [7:0] m_axi_rmem19_AWLEN;
  (* RS_HS = "m_axi_rmem19_AW.data" *)output m_axi_rmem19_AWLOCK;
  (* RS_HS = "m_axi_rmem19_AW.data" *)output [2:0] m_axi_rmem19_AWPROT;
  (* RS_HS = "m_axi_rmem19_AW.data" *)output [3:0] m_axi_rmem19_AWQOS;
  (* RS_HS = "m_axi_rmem19_AW.ready" *)input m_axi_rmem19_AWREADY;
  (* RS_HS = "m_axi_rmem19_AW.data" *)output [2:0] m_axi_rmem19_AWSIZE;
  (* RS_HS = "m_axi_rmem19_AW.valid" *)output m_axi_rmem19_AWVALID;
  (* RS_HS = "m_axi_rmem19_B.data" *)input [1:0] m_axi_rmem19_BID;
  (* RS_HS = "m_axi_rmem19_B.ready" *)output m_axi_rmem19_BREADY;
  (* RS_HS = "m_axi_rmem19_B.data" *)input [1:0] m_axi_rmem19_BRESP;
  (* RS_HS = "m_axi_rmem19_B.valid" *)input m_axi_rmem19_BVALID;
  (* RS_HS = "m_axi_rmem19_R.data" *)input [511:0] m_axi_rmem19_RDATA;
  (* RS_HS = "m_axi_rmem19_R.data" *)input [1:0] m_axi_rmem19_RID;
  (* RS_HS = "m_axi_rmem19_R.data" *)input m_axi_rmem19_RLAST;
  (* RS_HS = "m_axi_rmem19_R.ready" *)output m_axi_rmem19_RREADY;
  (* RS_HS = "m_axi_rmem19_R.data" *)input [1:0] m_axi_rmem19_RRESP;
  (* RS_HS = "m_axi_rmem19_R.valid" *)input m_axi_rmem19_RVALID;
  (* RS_HS = "m_axi_rmem19_W.data" *)output [511:0] m_axi_rmem19_WDATA;
  (* RS_HS = "m_axi_rmem19_W.data" *)output m_axi_rmem19_WLAST;
  (* RS_HS = "m_axi_rmem19_W.ready" *)input m_axi_rmem19_WREADY;
  (* RS_HS = "m_axi_rmem19_W.data" *)output [63:0] m_axi_rmem19_WSTRB;
  (* RS_HS = "m_axi_rmem19_W.valid" *)output m_axi_rmem19_WVALID;
  (* RS_HS = "m_axi_rmem20_AR.data" *)output [63:0] m_axi_rmem20_ARADDR;
  (* RS_HS = "m_axi_rmem20_AR.data" *)output [1:0] m_axi_rmem20_ARBURST;
  (* RS_HS = "m_axi_rmem20_AR.data" *)output [3:0] m_axi_rmem20_ARCACHE;
  (* RS_HS = "m_axi_rmem20_AR.data" *)output [1:0] m_axi_rmem20_ARID;
  (* RS_HS = "m_axi_rmem20_AR.data" *)output [7:0] m_axi_rmem20_ARLEN;
  (* RS_HS = "m_axi_rmem20_AR.data" *)output m_axi_rmem20_ARLOCK;
  (* RS_HS = "m_axi_rmem20_AR.data" *)output [2:0] m_axi_rmem20_ARPROT;
  (* RS_HS = "m_axi_rmem20_AR.data" *)output [3:0] m_axi_rmem20_ARQOS;
  (* RS_HS = "m_axi_rmem20_AR.ready" *)input m_axi_rmem20_ARREADY;
  (* RS_HS = "m_axi_rmem20_AR.data" *)output [2:0] m_axi_rmem20_ARSIZE;
  (* RS_HS = "m_axi_rmem20_AR.valid" *)output m_axi_rmem20_ARVALID;
  (* RS_HS = "m_axi_rmem20_AW.data" *)output [63:0] m_axi_rmem20_AWADDR;
  (* RS_HS = "m_axi_rmem20_AW.data" *)output [1:0] m_axi_rmem20_AWBURST;
  (* RS_HS = "m_axi_rmem20_AW.data" *)output [3:0] m_axi_rmem20_AWCACHE;
  (* RS_HS = "m_axi_rmem20_AW.data" *)output [1:0] m_axi_rmem20_AWID;
  (* RS_HS = "m_axi_rmem20_AW.data" *)output [7:0] m_axi_rmem20_AWLEN;
  (* RS_HS = "m_axi_rmem20_AW.data" *)output m_axi_rmem20_AWLOCK;
  (* RS_HS = "m_axi_rmem20_AW.data" *)output [2:0] m_axi_rmem20_AWPROT;
  (* RS_HS = "m_axi_rmem20_AW.data" *)output [3:0] m_axi_rmem20_AWQOS;
  (* RS_HS = "m_axi_rmem20_AW.ready" *)input m_axi_rmem20_AWREADY;
  (* RS_HS = "m_axi_rmem20_AW.data" *)output [2:0] m_axi_rmem20_AWSIZE;
  (* RS_HS = "m_axi_rmem20_AW.valid" *)output m_axi_rmem20_AWVALID;
  (* RS_HS = "m_axi_rmem20_B.data" *)input [1:0] m_axi_rmem20_BID;
  (* RS_HS = "m_axi_rmem20_B.ready" *)output m_axi_rmem20_BREADY;
  (* RS_HS = "m_axi_rmem20_B.data" *)input [1:0] m_axi_rmem20_BRESP;
  (* RS_HS = "m_axi_rmem20_B.valid" *)input m_axi_rmem20_BVALID;
  (* RS_HS = "m_axi_rmem20_R.data" *)input [511:0] m_axi_rmem20_RDATA;
  (* RS_HS = "m_axi_rmem20_R.data" *)input [1:0] m_axi_rmem20_RID;
  (* RS_HS = "m_axi_rmem20_R.data" *)input m_axi_rmem20_RLAST;
  (* RS_HS = "m_axi_rmem20_R.ready" *)output m_axi_rmem20_RREADY;
  (* RS_HS = "m_axi_rmem20_R.data" *)input [1:0] m_axi_rmem20_RRESP;
  (* RS_HS = "m_axi_rmem20_R.valid" *)input m_axi_rmem20_RVALID;
  (* RS_HS = "m_axi_rmem20_W.data" *)output [511:0] m_axi_rmem20_WDATA;
  (* RS_HS = "m_axi_rmem20_W.data" *)output m_axi_rmem20_WLAST;
  (* RS_HS = "m_axi_rmem20_W.ready" *)input m_axi_rmem20_WREADY;
  (* RS_HS = "m_axi_rmem20_W.data" *)output [63:0] m_axi_rmem20_WSTRB;
  (* RS_HS = "m_axi_rmem20_W.valid" *)output m_axi_rmem20_WVALID;
  (* RS_HS = "m_axi_rmem21_AR.data" *)output [63:0] m_axi_rmem21_ARADDR;
  (* RS_HS = "m_axi_rmem21_AR.data" *)output [1:0] m_axi_rmem21_ARBURST;
  (* RS_HS = "m_axi_rmem21_AR.data" *)output [3:0] m_axi_rmem21_ARCACHE;
  (* RS_HS = "m_axi_rmem21_AR.data" *)output [1:0] m_axi_rmem21_ARID;
  (* RS_HS = "m_axi_rmem21_AR.data" *)output [7:0] m_axi_rmem21_ARLEN;
  (* RS_HS = "m_axi_rmem21_AR.data" *)output m_axi_rmem21_ARLOCK;
  (* RS_HS = "m_axi_rmem21_AR.data" *)output [2:0] m_axi_rmem21_ARPROT;
  (* RS_HS = "m_axi_rmem21_AR.data" *)output [3:0] m_axi_rmem21_ARQOS;
  (* RS_HS = "m_axi_rmem21_AR.ready" *)input m_axi_rmem21_ARREADY;
  (* RS_HS = "m_axi_rmem21_AR.data" *)output [2:0] m_axi_rmem21_ARSIZE;
  (* RS_HS = "m_axi_rmem21_AR.valid" *)output m_axi_rmem21_ARVALID;
  (* RS_HS = "m_axi_rmem21_AW.data" *)output [63:0] m_axi_rmem21_AWADDR;
  (* RS_HS = "m_axi_rmem21_AW.data" *)output [1:0] m_axi_rmem21_AWBURST;
  (* RS_HS = "m_axi_rmem21_AW.data" *)output [3:0] m_axi_rmem21_AWCACHE;
  (* RS_HS = "m_axi_rmem21_AW.data" *)output [1:0] m_axi_rmem21_AWID;
  (* RS_HS = "m_axi_rmem21_AW.data" *)output [7:0] m_axi_rmem21_AWLEN;
  (* RS_HS = "m_axi_rmem21_AW.data" *)output m_axi_rmem21_AWLOCK;
  (* RS_HS = "m_axi_rmem21_AW.data" *)output [2:0] m_axi_rmem21_AWPROT;
  (* RS_HS = "m_axi_rmem21_AW.data" *)output [3:0] m_axi_rmem21_AWQOS;
  (* RS_HS = "m_axi_rmem21_AW.ready" *)input m_axi_rmem21_AWREADY;
  (* RS_HS = "m_axi_rmem21_AW.data" *)output [2:0] m_axi_rmem21_AWSIZE;
  (* RS_HS = "m_axi_rmem21_AW.valid" *)output m_axi_rmem21_AWVALID;
  (* RS_HS = "m_axi_rmem21_B.data" *)input [1:0] m_axi_rmem21_BID;
  (* RS_HS = "m_axi_rmem21_B.ready" *)output m_axi_rmem21_BREADY;
  (* RS_HS = "m_axi_rmem21_B.data" *)input [1:0] m_axi_rmem21_BRESP;
  (* RS_HS = "m_axi_rmem21_B.valid" *)input m_axi_rmem21_BVALID;
  (* RS_HS = "m_axi_rmem21_R.data" *)input [511:0] m_axi_rmem21_RDATA;
  (* RS_HS = "m_axi_rmem21_R.data" *)input [1:0] m_axi_rmem21_RID;
  (* RS_HS = "m_axi_rmem21_R.data" *)input m_axi_rmem21_RLAST;
  (* RS_HS = "m_axi_rmem21_R.ready" *)output m_axi_rmem21_RREADY;
  (* RS_HS = "m_axi_rmem21_R.data" *)input [1:0] m_axi_rmem21_RRESP;
  (* RS_HS = "m_axi_rmem21_R.valid" *)input m_axi_rmem21_RVALID;
  (* RS_HS = "m_axi_rmem21_W.data" *)output [511:0] m_axi_rmem21_WDATA;
  (* RS_HS = "m_axi_rmem21_W.data" *)output m_axi_rmem21_WLAST;
  (* RS_HS = "m_axi_rmem21_W.ready" *)input m_axi_rmem21_WREADY;
  (* RS_HS = "m_axi_rmem21_W.data" *)output [63:0] m_axi_rmem21_WSTRB;
  (* RS_HS = "m_axi_rmem21_W.valid" *)output m_axi_rmem21_WVALID;
  (* RS_HS = "m_axi_rmem22_AR.data" *)output [63:0] m_axi_rmem22_ARADDR;
  (* RS_HS = "m_axi_rmem22_AR.data" *)output [1:0] m_axi_rmem22_ARBURST;
  (* RS_HS = "m_axi_rmem22_AR.data" *)output [3:0] m_axi_rmem22_ARCACHE;
  (* RS_HS = "m_axi_rmem22_AR.data" *)output [1:0] m_axi_rmem22_ARID;
  (* RS_HS = "m_axi_rmem22_AR.data" *)output [7:0] m_axi_rmem22_ARLEN;
  (* RS_HS = "m_axi_rmem22_AR.data" *)output m_axi_rmem22_ARLOCK;
  (* RS_HS = "m_axi_rmem22_AR.data" *)output [2:0] m_axi_rmem22_ARPROT;
  (* RS_HS = "m_axi_rmem22_AR.data" *)output [3:0] m_axi_rmem22_ARQOS;
  (* RS_HS = "m_axi_rmem22_AR.ready" *)input m_axi_rmem22_ARREADY;
  (* RS_HS = "m_axi_rmem22_AR.data" *)output [2:0] m_axi_rmem22_ARSIZE;
  (* RS_HS = "m_axi_rmem22_AR.valid" *)output m_axi_rmem22_ARVALID;
  (* RS_HS = "m_axi_rmem22_AW.data" *)output [63:0] m_axi_rmem22_AWADDR;
  (* RS_HS = "m_axi_rmem22_AW.data" *)output [1:0] m_axi_rmem22_AWBURST;
  (* RS_HS = "m_axi_rmem22_AW.data" *)output [3:0] m_axi_rmem22_AWCACHE;
  (* RS_HS = "m_axi_rmem22_AW.data" *)output [1:0] m_axi_rmem22_AWID;
  (* RS_HS = "m_axi_rmem22_AW.data" *)output [7:0] m_axi_rmem22_AWLEN;
  (* RS_HS = "m_axi_rmem22_AW.data" *)output m_axi_rmem22_AWLOCK;
  (* RS_HS = "m_axi_rmem22_AW.data" *)output [2:0] m_axi_rmem22_AWPROT;
  (* RS_HS = "m_axi_rmem22_AW.data" *)output [3:0] m_axi_rmem22_AWQOS;
  (* RS_HS = "m_axi_rmem22_AW.ready" *)input m_axi_rmem22_AWREADY;
  (* RS_HS = "m_axi_rmem22_AW.data" *)output [2:0] m_axi_rmem22_AWSIZE;
  (* RS_HS = "m_axi_rmem22_AW.valid" *)output m_axi_rmem22_AWVALID;
  (* RS_HS = "m_axi_rmem22_B.data" *)input [1:0] m_axi_rmem22_BID;
  (* RS_HS = "m_axi_rmem22_B.ready" *)output m_axi_rmem22_BREADY;
  (* RS_HS = "m_axi_rmem22_B.data" *)input [1:0] m_axi_rmem22_BRESP;
  (* RS_HS = "m_axi_rmem22_B.valid" *)input m_axi_rmem22_BVALID;
  (* RS_HS = "m_axi_rmem22_R.data" *)input [511:0] m_axi_rmem22_RDATA;
  (* RS_HS = "m_axi_rmem22_R.data" *)input [1:0] m_axi_rmem22_RID;
  (* RS_HS = "m_axi_rmem22_R.data" *)input m_axi_rmem22_RLAST;
  (* RS_HS = "m_axi_rmem22_R.ready" *)output m_axi_rmem22_RREADY;
  (* RS_HS = "m_axi_rmem22_R.data" *)input [1:0] m_axi_rmem22_RRESP;
  (* RS_HS = "m_axi_rmem22_R.valid" *)input m_axi_rmem22_RVALID;
  (* RS_HS = "m_axi_rmem22_W.data" *)output [511:0] m_axi_rmem22_WDATA;
  (* RS_HS = "m_axi_rmem22_W.data" *)output m_axi_rmem22_WLAST;
  (* RS_HS = "m_axi_rmem22_W.ready" *)input m_axi_rmem22_WREADY;
  (* RS_HS = "m_axi_rmem22_W.data" *)output [63:0] m_axi_rmem22_WSTRB;
  (* RS_HS = "m_axi_rmem22_W.valid" *)output m_axi_rmem22_WVALID;
  (* RS_HS = "m_axi_rmem23_AR.data" *)output [63:0] m_axi_rmem23_ARADDR;
  (* RS_HS = "m_axi_rmem23_AR.data" *)output [1:0] m_axi_rmem23_ARBURST;
  (* RS_HS = "m_axi_rmem23_AR.data" *)output [3:0] m_axi_rmem23_ARCACHE;
  (* RS_HS = "m_axi_rmem23_AR.data" *)output [1:0] m_axi_rmem23_ARID;
  (* RS_HS = "m_axi_rmem23_AR.data" *)output [7:0] m_axi_rmem23_ARLEN;
  (* RS_HS = "m_axi_rmem23_AR.data" *)output m_axi_rmem23_ARLOCK;
  (* RS_HS = "m_axi_rmem23_AR.data" *)output [2:0] m_axi_rmem23_ARPROT;
  (* RS_HS = "m_axi_rmem23_AR.data" *)output [3:0] m_axi_rmem23_ARQOS;
  (* RS_HS = "m_axi_rmem23_AR.ready" *)input m_axi_rmem23_ARREADY;
  (* RS_HS = "m_axi_rmem23_AR.data" *)output [2:0] m_axi_rmem23_ARSIZE;
  (* RS_HS = "m_axi_rmem23_AR.valid" *)output m_axi_rmem23_ARVALID;
  (* RS_HS = "m_axi_rmem23_AW.data" *)output [63:0] m_axi_rmem23_AWADDR;
  (* RS_HS = "m_axi_rmem23_AW.data" *)output [1:0] m_axi_rmem23_AWBURST;
  (* RS_HS = "m_axi_rmem23_AW.data" *)output [3:0] m_axi_rmem23_AWCACHE;
  (* RS_HS = "m_axi_rmem23_AW.data" *)output [1:0] m_axi_rmem23_AWID;
  (* RS_HS = "m_axi_rmem23_AW.data" *)output [7:0] m_axi_rmem23_AWLEN;
  (* RS_HS = "m_axi_rmem23_AW.data" *)output m_axi_rmem23_AWLOCK;
  (* RS_HS = "m_axi_rmem23_AW.data" *)output [2:0] m_axi_rmem23_AWPROT;
  (* RS_HS = "m_axi_rmem23_AW.data" *)output [3:0] m_axi_rmem23_AWQOS;
  (* RS_HS = "m_axi_rmem23_AW.ready" *)input m_axi_rmem23_AWREADY;
  (* RS_HS = "m_axi_rmem23_AW.data" *)output [2:0] m_axi_rmem23_AWSIZE;
  (* RS_HS = "m_axi_rmem23_AW.valid" *)output m_axi_rmem23_AWVALID;
  (* RS_HS = "m_axi_rmem23_B.data" *)input [1:0] m_axi_rmem23_BID;
  (* RS_HS = "m_axi_rmem23_B.ready" *)output m_axi_rmem23_BREADY;
  (* RS_HS = "m_axi_rmem23_B.data" *)input [1:0] m_axi_rmem23_BRESP;
  (* RS_HS = "m_axi_rmem23_B.valid" *)input m_axi_rmem23_BVALID;
  (* RS_HS = "m_axi_rmem23_R.data" *)input [511:0] m_axi_rmem23_RDATA;
  (* RS_HS = "m_axi_rmem23_R.data" *)input [1:0] m_axi_rmem23_RID;
  (* RS_HS = "m_axi_rmem23_R.data" *)input m_axi_rmem23_RLAST;
  (* RS_HS = "m_axi_rmem23_R.ready" *)output m_axi_rmem23_RREADY;
  (* RS_HS = "m_axi_rmem23_R.data" *)input [1:0] m_axi_rmem23_RRESP;
  (* RS_HS = "m_axi_rmem23_R.valid" *)input m_axi_rmem23_RVALID;
  (* RS_HS = "m_axi_rmem23_W.data" *)output [511:0] m_axi_rmem23_WDATA;
  (* RS_HS = "m_axi_rmem23_W.data" *)output m_axi_rmem23_WLAST;
  (* RS_HS = "m_axi_rmem23_W.ready" *)input m_axi_rmem23_WREADY;
  (* RS_HS = "m_axi_rmem23_W.data" *)output [63:0] m_axi_rmem23_WSTRB;
  (* RS_HS = "m_axi_rmem23_W.valid" *)output m_axi_rmem23_WVALID;
  (* RS_HS = "m_axi_rmem24_AR.data" *)output [63:0] m_axi_rmem24_ARADDR;
  (* RS_HS = "m_axi_rmem24_AR.data" *)output [1:0] m_axi_rmem24_ARBURST;
  (* RS_HS = "m_axi_rmem24_AR.data" *)output [3:0] m_axi_rmem24_ARCACHE;
  (* RS_HS = "m_axi_rmem24_AR.data" *)output [1:0] m_axi_rmem24_ARID;
  (* RS_HS = "m_axi_rmem24_AR.data" *)output [7:0] m_axi_rmem24_ARLEN;
  (* RS_HS = "m_axi_rmem24_AR.data" *)output m_axi_rmem24_ARLOCK;
  (* RS_HS = "m_axi_rmem24_AR.data" *)output [2:0] m_axi_rmem24_ARPROT;
  (* RS_HS = "m_axi_rmem24_AR.data" *)output [3:0] m_axi_rmem24_ARQOS;
  (* RS_HS = "m_axi_rmem24_AR.ready" *)input m_axi_rmem24_ARREADY;
  (* RS_HS = "m_axi_rmem24_AR.data" *)output [2:0] m_axi_rmem24_ARSIZE;
  (* RS_HS = "m_axi_rmem24_AR.valid" *)output m_axi_rmem24_ARVALID;
  (* RS_HS = "m_axi_rmem24_AW.data" *)output [63:0] m_axi_rmem24_AWADDR;
  (* RS_HS = "m_axi_rmem24_AW.data" *)output [1:0] m_axi_rmem24_AWBURST;
  (* RS_HS = "m_axi_rmem24_AW.data" *)output [3:0] m_axi_rmem24_AWCACHE;
  (* RS_HS = "m_axi_rmem24_AW.data" *)output [1:0] m_axi_rmem24_AWID;
  (* RS_HS = "m_axi_rmem24_AW.data" *)output [7:0] m_axi_rmem24_AWLEN;
  (* RS_HS = "m_axi_rmem24_AW.data" *)output m_axi_rmem24_AWLOCK;
  (* RS_HS = "m_axi_rmem24_AW.data" *)output [2:0] m_axi_rmem24_AWPROT;
  (* RS_HS = "m_axi_rmem24_AW.data" *)output [3:0] m_axi_rmem24_AWQOS;
  (* RS_HS = "m_axi_rmem24_AW.ready" *)input m_axi_rmem24_AWREADY;
  (* RS_HS = "m_axi_rmem24_AW.data" *)output [2:0] m_axi_rmem24_AWSIZE;
  (* RS_HS = "m_axi_rmem24_AW.valid" *)output m_axi_rmem24_AWVALID;
  (* RS_HS = "m_axi_rmem24_B.data" *)input [1:0] m_axi_rmem24_BID;
  (* RS_HS = "m_axi_rmem24_B.ready" *)output m_axi_rmem24_BREADY;
  (* RS_HS = "m_axi_rmem24_B.data" *)input [1:0] m_axi_rmem24_BRESP;
  (* RS_HS = "m_axi_rmem24_B.valid" *)input m_axi_rmem24_BVALID;
  (* RS_HS = "m_axi_rmem24_R.data" *)input [511:0] m_axi_rmem24_RDATA;
  (* RS_HS = "m_axi_rmem24_R.data" *)input [1:0] m_axi_rmem24_RID;
  (* RS_HS = "m_axi_rmem24_R.data" *)input m_axi_rmem24_RLAST;
  (* RS_HS = "m_axi_rmem24_R.ready" *)output m_axi_rmem24_RREADY;
  (* RS_HS = "m_axi_rmem24_R.data" *)input [1:0] m_axi_rmem24_RRESP;
  (* RS_HS = "m_axi_rmem24_R.valid" *)input m_axi_rmem24_RVALID;
  (* RS_HS = "m_axi_rmem24_W.data" *)output [511:0] m_axi_rmem24_WDATA;
  (* RS_HS = "m_axi_rmem24_W.data" *)output m_axi_rmem24_WLAST;
  (* RS_HS = "m_axi_rmem24_W.ready" *)input m_axi_rmem24_WREADY;
  (* RS_HS = "m_axi_rmem24_W.data" *)output [63:0] m_axi_rmem24_WSTRB;
  (* RS_HS = "m_axi_rmem24_W.valid" *)output m_axi_rmem24_WVALID;
  (* RS_HS = "m_axi_rmem25_AR.data" *)output [63:0] m_axi_rmem25_ARADDR;
  (* RS_HS = "m_axi_rmem25_AR.data" *)output [1:0] m_axi_rmem25_ARBURST;
  (* RS_HS = "m_axi_rmem25_AR.data" *)output [3:0] m_axi_rmem25_ARCACHE;
  (* RS_HS = "m_axi_rmem25_AR.data" *)output [1:0] m_axi_rmem25_ARID;
  (* RS_HS = "m_axi_rmem25_AR.data" *)output [7:0] m_axi_rmem25_ARLEN;
  (* RS_HS = "m_axi_rmem25_AR.data" *)output m_axi_rmem25_ARLOCK;
  (* RS_HS = "m_axi_rmem25_AR.data" *)output [2:0] m_axi_rmem25_ARPROT;
  (* RS_HS = "m_axi_rmem25_AR.data" *)output [3:0] m_axi_rmem25_ARQOS;
  (* RS_HS = "m_axi_rmem25_AR.ready" *)input m_axi_rmem25_ARREADY;
  (* RS_HS = "m_axi_rmem25_AR.data" *)output [2:0] m_axi_rmem25_ARSIZE;
  (* RS_HS = "m_axi_rmem25_AR.valid" *)output m_axi_rmem25_ARVALID;
  (* RS_HS = "m_axi_rmem25_AW.data" *)output [63:0] m_axi_rmem25_AWADDR;
  (* RS_HS = "m_axi_rmem25_AW.data" *)output [1:0] m_axi_rmem25_AWBURST;
  (* RS_HS = "m_axi_rmem25_AW.data" *)output [3:0] m_axi_rmem25_AWCACHE;
  (* RS_HS = "m_axi_rmem25_AW.data" *)output [1:0] m_axi_rmem25_AWID;
  (* RS_HS = "m_axi_rmem25_AW.data" *)output [7:0] m_axi_rmem25_AWLEN;
  (* RS_HS = "m_axi_rmem25_AW.data" *)output m_axi_rmem25_AWLOCK;
  (* RS_HS = "m_axi_rmem25_AW.data" *)output [2:0] m_axi_rmem25_AWPROT;
  (* RS_HS = "m_axi_rmem25_AW.data" *)output [3:0] m_axi_rmem25_AWQOS;
  (* RS_HS = "m_axi_rmem25_AW.ready" *)input m_axi_rmem25_AWREADY;
  (* RS_HS = "m_axi_rmem25_AW.data" *)output [2:0] m_axi_rmem25_AWSIZE;
  (* RS_HS = "m_axi_rmem25_AW.valid" *)output m_axi_rmem25_AWVALID;
  (* RS_HS = "m_axi_rmem25_B.data" *)input [1:0] m_axi_rmem25_BID;
  (* RS_HS = "m_axi_rmem25_B.ready" *)output m_axi_rmem25_BREADY;
  (* RS_HS = "m_axi_rmem25_B.data" *)input [1:0] m_axi_rmem25_BRESP;
  (* RS_HS = "m_axi_rmem25_B.valid" *)input m_axi_rmem25_BVALID;
  (* RS_HS = "m_axi_rmem25_R.data" *)input [511:0] m_axi_rmem25_RDATA;
  (* RS_HS = "m_axi_rmem25_R.data" *)input [1:0] m_axi_rmem25_RID;
  (* RS_HS = "m_axi_rmem25_R.data" *)input m_axi_rmem25_RLAST;
  (* RS_HS = "m_axi_rmem25_R.ready" *)output m_axi_rmem25_RREADY;
  (* RS_HS = "m_axi_rmem25_R.data" *)input [1:0] m_axi_rmem25_RRESP;
  (* RS_HS = "m_axi_rmem25_R.valid" *)input m_axi_rmem25_RVALID;
  (* RS_HS = "m_axi_rmem25_W.data" *)output [511:0] m_axi_rmem25_WDATA;
  (* RS_HS = "m_axi_rmem25_W.data" *)output m_axi_rmem25_WLAST;
  (* RS_HS = "m_axi_rmem25_W.ready" *)input m_axi_rmem25_WREADY;
  (* RS_HS = "m_axi_rmem25_W.data" *)output [63:0] m_axi_rmem25_WSTRB;
  (* RS_HS = "m_axi_rmem25_W.valid" *)output m_axi_rmem25_WVALID;
  (* RS_HS = "m_axi_rmem26_AR.data" *)output [63:0] m_axi_rmem26_ARADDR;
  (* RS_HS = "m_axi_rmem26_AR.data" *)output [1:0] m_axi_rmem26_ARBURST;
  (* RS_HS = "m_axi_rmem26_AR.data" *)output [3:0] m_axi_rmem26_ARCACHE;
  (* RS_HS = "m_axi_rmem26_AR.data" *)output [1:0] m_axi_rmem26_ARID;
  (* RS_HS = "m_axi_rmem26_AR.data" *)output [7:0] m_axi_rmem26_ARLEN;
  (* RS_HS = "m_axi_rmem26_AR.data" *)output m_axi_rmem26_ARLOCK;
  (* RS_HS = "m_axi_rmem26_AR.data" *)output [2:0] m_axi_rmem26_ARPROT;
  (* RS_HS = "m_axi_rmem26_AR.data" *)output [3:0] m_axi_rmem26_ARQOS;
  (* RS_HS = "m_axi_rmem26_AR.ready" *)input m_axi_rmem26_ARREADY;
  (* RS_HS = "m_axi_rmem26_AR.data" *)output [2:0] m_axi_rmem26_ARSIZE;
  (* RS_HS = "m_axi_rmem26_AR.valid" *)output m_axi_rmem26_ARVALID;
  (* RS_HS = "m_axi_rmem26_AW.data" *)output [63:0] m_axi_rmem26_AWADDR;
  (* RS_HS = "m_axi_rmem26_AW.data" *)output [1:0] m_axi_rmem26_AWBURST;
  (* RS_HS = "m_axi_rmem26_AW.data" *)output [3:0] m_axi_rmem26_AWCACHE;
  (* RS_HS = "m_axi_rmem26_AW.data" *)output [1:0] m_axi_rmem26_AWID;
  (* RS_HS = "m_axi_rmem26_AW.data" *)output [7:0] m_axi_rmem26_AWLEN;
  (* RS_HS = "m_axi_rmem26_AW.data" *)output m_axi_rmem26_AWLOCK;
  (* RS_HS = "m_axi_rmem26_AW.data" *)output [2:0] m_axi_rmem26_AWPROT;
  (* RS_HS = "m_axi_rmem26_AW.data" *)output [3:0] m_axi_rmem26_AWQOS;
  (* RS_HS = "m_axi_rmem26_AW.ready" *)input m_axi_rmem26_AWREADY;
  (* RS_HS = "m_axi_rmem26_AW.data" *)output [2:0] m_axi_rmem26_AWSIZE;
  (* RS_HS = "m_axi_rmem26_AW.valid" *)output m_axi_rmem26_AWVALID;
  (* RS_HS = "m_axi_rmem26_B.data" *)input [1:0] m_axi_rmem26_BID;
  (* RS_HS = "m_axi_rmem26_B.ready" *)output m_axi_rmem26_BREADY;
  (* RS_HS = "m_axi_rmem26_B.data" *)input [1:0] m_axi_rmem26_BRESP;
  (* RS_HS = "m_axi_rmem26_B.valid" *)input m_axi_rmem26_BVALID;
  (* RS_HS = "m_axi_rmem26_R.data" *)input [511:0] m_axi_rmem26_RDATA;
  (* RS_HS = "m_axi_rmem26_R.data" *)input [1:0] m_axi_rmem26_RID;
  (* RS_HS = "m_axi_rmem26_R.data" *)input m_axi_rmem26_RLAST;
  (* RS_HS = "m_axi_rmem26_R.ready" *)output m_axi_rmem26_RREADY;
  (* RS_HS = "m_axi_rmem26_R.data" *)input [1:0] m_axi_rmem26_RRESP;
  (* RS_HS = "m_axi_rmem26_R.valid" *)input m_axi_rmem26_RVALID;
  (* RS_HS = "m_axi_rmem26_W.data" *)output [511:0] m_axi_rmem26_WDATA;
  (* RS_HS = "m_axi_rmem26_W.data" *)output m_axi_rmem26_WLAST;
  (* RS_HS = "m_axi_rmem26_W.ready" *)input m_axi_rmem26_WREADY;
  (* RS_HS = "m_axi_rmem26_W.data" *)output [63:0] m_axi_rmem26_WSTRB;
  (* RS_HS = "m_axi_rmem26_W.valid" *)output m_axi_rmem26_WVALID;
  (* RS_HS = "m_axi_rmem27_AR.data" *)output [63:0] m_axi_rmem27_ARADDR;
  (* RS_HS = "m_axi_rmem27_AR.data" *)output [1:0] m_axi_rmem27_ARBURST;
  (* RS_HS = "m_axi_rmem27_AR.data" *)output [3:0] m_axi_rmem27_ARCACHE;
  (* RS_HS = "m_axi_rmem27_AR.data" *)output [1:0] m_axi_rmem27_ARID;
  (* RS_HS = "m_axi_rmem27_AR.data" *)output [7:0] m_axi_rmem27_ARLEN;
  (* RS_HS = "m_axi_rmem27_AR.data" *)output m_axi_rmem27_ARLOCK;
  (* RS_HS = "m_axi_rmem27_AR.data" *)output [2:0] m_axi_rmem27_ARPROT;
  (* RS_HS = "m_axi_rmem27_AR.data" *)output [3:0] m_axi_rmem27_ARQOS;
  (* RS_HS = "m_axi_rmem27_AR.ready" *)input m_axi_rmem27_ARREADY;
  (* RS_HS = "m_axi_rmem27_AR.data" *)output [2:0] m_axi_rmem27_ARSIZE;
  (* RS_HS = "m_axi_rmem27_AR.valid" *)output m_axi_rmem27_ARVALID;
  (* RS_HS = "m_axi_rmem27_AW.data" *)output [63:0] m_axi_rmem27_AWADDR;
  (* RS_HS = "m_axi_rmem27_AW.data" *)output [1:0] m_axi_rmem27_AWBURST;
  (* RS_HS = "m_axi_rmem27_AW.data" *)output [3:0] m_axi_rmem27_AWCACHE;
  (* RS_HS = "m_axi_rmem27_AW.data" *)output [1:0] m_axi_rmem27_AWID;
  (* RS_HS = "m_axi_rmem27_AW.data" *)output [7:0] m_axi_rmem27_AWLEN;
  (* RS_HS = "m_axi_rmem27_AW.data" *)output m_axi_rmem27_AWLOCK;
  (* RS_HS = "m_axi_rmem27_AW.data" *)output [2:0] m_axi_rmem27_AWPROT;
  (* RS_HS = "m_axi_rmem27_AW.data" *)output [3:0] m_axi_rmem27_AWQOS;
  (* RS_HS = "m_axi_rmem27_AW.ready" *)input m_axi_rmem27_AWREADY;
  (* RS_HS = "m_axi_rmem27_AW.data" *)output [2:0] m_axi_rmem27_AWSIZE;
  (* RS_HS = "m_axi_rmem27_AW.valid" *)output m_axi_rmem27_AWVALID;
  (* RS_HS = "m_axi_rmem27_B.data" *)input [1:0] m_axi_rmem27_BID;
  (* RS_HS = "m_axi_rmem27_B.ready" *)output m_axi_rmem27_BREADY;
  (* RS_HS = "m_axi_rmem27_B.data" *)input [1:0] m_axi_rmem27_BRESP;
  (* RS_HS = "m_axi_rmem27_B.valid" *)input m_axi_rmem27_BVALID;
  (* RS_HS = "m_axi_rmem27_R.data" *)input [511:0] m_axi_rmem27_RDATA;
  (* RS_HS = "m_axi_rmem27_R.data" *)input [1:0] m_axi_rmem27_RID;
  (* RS_HS = "m_axi_rmem27_R.data" *)input m_axi_rmem27_RLAST;
  (* RS_HS = "m_axi_rmem27_R.ready" *)output m_axi_rmem27_RREADY;
  (* RS_HS = "m_axi_rmem27_R.data" *)input [1:0] m_axi_rmem27_RRESP;
  (* RS_HS = "m_axi_rmem27_R.valid" *)input m_axi_rmem27_RVALID;
  (* RS_HS = "m_axi_rmem27_W.data" *)output [511:0] m_axi_rmem27_WDATA;
  (* RS_HS = "m_axi_rmem27_W.data" *)output m_axi_rmem27_WLAST;
  (* RS_HS = "m_axi_rmem27_W.ready" *)input m_axi_rmem27_WREADY;
  (* RS_HS = "m_axi_rmem27_W.data" *)output [63:0] m_axi_rmem27_WSTRB;
  (* RS_HS = "m_axi_rmem27_W.valid" *)output m_axi_rmem27_WVALID;
  wire ap_start;
  wire [63:0] rmem0;
  wire [63:0] rmem1;
  wire [63:0] rmem2;
  wire [63:0] rmem3;
  wire [63:0] rmem4;
  wire [63:0] rmem5;
  wire [63:0] rmem6;
  wire [63:0] rmem7;
  wire [63:0] rmem8;
  wire [63:0] rmem9;
  wire [63:0] rmem10;
  wire [63:0] rmem11;
  wire [63:0] rmem12;
  wire [63:0] rmem13;
  wire [63:0] rmem14;
  wire [63:0] rmem15;
  wire [63:0] rmem16;
  wire [63:0] rmem17;
  wire [63:0] rmem18;
  wire [63:0] rmem19;
  wire [63:0] rmem20;
  wire [63:0] rmem21;
  wire [63:0] rmem22;
  wire [63:0] rmem23;
  wire [63:0] rmem24;
  wire [63:0] rmem25;
  wire [63:0] rmem26;
  wire [63:0] rmem27;
  wire [63:0] n;
  wire [512:0] qr0_vadd_bw__dout;
  wire qr0_vadd_bw__empty_n;
  wire qr0_vadd_bw__read;
  wire [512:0] qr0_vadd_bw__din;
  wire qr0_vadd_bw__full_n;
  wire qr0_vadd_bw__write;
  wire [512:0] qr10_vadd_bw__dout;
  wire qr10_vadd_bw__empty_n;
  wire qr10_vadd_bw__read;
  wire [512:0] qr10_vadd_bw__din;
  wire qr10_vadd_bw__full_n;
  wire qr10_vadd_bw__write;
  wire [512:0] qr11_vadd_bw__dout;
  wire qr11_vadd_bw__empty_n;
  wire qr11_vadd_bw__read;
  wire [512:0] qr11_vadd_bw__din;
  wire qr11_vadd_bw__full_n;
  wire qr11_vadd_bw__write;
  wire [512:0] qr12_vadd_bw__dout;
  wire qr12_vadd_bw__empty_n;
  wire qr12_vadd_bw__read;
  wire [512:0] qr12_vadd_bw__din;
  wire qr12_vadd_bw__full_n;
  wire qr12_vadd_bw__write;
  wire [512:0] qr13_vadd_bw__dout;
  wire qr13_vadd_bw__empty_n;
  wire qr13_vadd_bw__read;
  wire [512:0] qr13_vadd_bw__din;
  wire qr13_vadd_bw__full_n;
  wire qr13_vadd_bw__write;
  wire [512:0] qr14_vadd_bw__dout;
  wire qr14_vadd_bw__empty_n;
  wire qr14_vadd_bw__read;
  wire [512:0] qr14_vadd_bw__din;
  wire qr14_vadd_bw__full_n;
  wire qr14_vadd_bw__write;
  wire [512:0] qr15_vadd_bw__dout;
  wire qr15_vadd_bw__empty_n;
  wire qr15_vadd_bw__read;
  wire [512:0] qr15_vadd_bw__din;
  wire qr15_vadd_bw__full_n;
  wire qr15_vadd_bw__write;
  wire [512:0] qr16_vadd_bw__dout;
  wire qr16_vadd_bw__empty_n;
  wire qr16_vadd_bw__read;
  wire [512:0] qr16_vadd_bw__din;
  wire qr16_vadd_bw__full_n;
  wire qr16_vadd_bw__write;
  wire [512:0] qr17_vadd_bw__dout;
  wire qr17_vadd_bw__empty_n;
  wire qr17_vadd_bw__read;
  wire [512:0] qr17_vadd_bw__din;
  wire qr17_vadd_bw__full_n;
  wire qr17_vadd_bw__write;
  wire [512:0] qr18_vadd_bw__dout;
  wire qr18_vadd_bw__empty_n;
  wire qr18_vadd_bw__read;
  wire [512:0] qr18_vadd_bw__din;
  wire qr18_vadd_bw__full_n;
  wire qr18_vadd_bw__write;
  wire [512:0] qr19_vadd_bw__dout;
  wire qr19_vadd_bw__empty_n;
  wire qr19_vadd_bw__read;
  wire [512:0] qr19_vadd_bw__din;
  wire qr19_vadd_bw__full_n;
  wire qr19_vadd_bw__write;
  wire [512:0] qr1_vadd_bw__dout;
  wire qr1_vadd_bw__empty_n;
  wire qr1_vadd_bw__read;
  wire [512:0] qr1_vadd_bw__din;
  wire qr1_vadd_bw__full_n;
  wire qr1_vadd_bw__write;
  wire [512:0] qr20_vadd_bw__dout;
  wire qr20_vadd_bw__empty_n;
  wire qr20_vadd_bw__read;
  wire [512:0] qr20_vadd_bw__din;
  wire qr20_vadd_bw__full_n;
  wire qr20_vadd_bw__write;
  wire [512:0] qr21_vadd_bw__dout;
  wire qr21_vadd_bw__empty_n;
  wire qr21_vadd_bw__read;
  wire [512:0] qr21_vadd_bw__din;
  wire qr21_vadd_bw__full_n;
  wire qr21_vadd_bw__write;
  wire [512:0] qr22_vadd_bw__dout;
  wire qr22_vadd_bw__empty_n;
  wire qr22_vadd_bw__read;
  wire [512:0] qr22_vadd_bw__din;
  wire qr22_vadd_bw__full_n;
  wire qr22_vadd_bw__write;
  wire [512:0] qr23_vadd_bw__dout;
  wire qr23_vadd_bw__empty_n;
  wire qr23_vadd_bw__read;
  wire [512:0] qr23_vadd_bw__din;
  wire qr23_vadd_bw__full_n;
  wire qr23_vadd_bw__write;
  wire [512:0] qr24_vadd_bw__dout;
  wire qr24_vadd_bw__empty_n;
  wire qr24_vadd_bw__read;
  wire [512:0] qr24_vadd_bw__din;
  wire qr24_vadd_bw__full_n;
  wire qr24_vadd_bw__write;
  wire [512:0] qr25_vadd_bw__dout;
  wire qr25_vadd_bw__empty_n;
  wire qr25_vadd_bw__read;
  wire [512:0] qr25_vadd_bw__din;
  wire qr25_vadd_bw__full_n;
  wire qr25_vadd_bw__write;
  wire [512:0] qr26_vadd_bw__dout;
  wire qr26_vadd_bw__empty_n;
  wire qr26_vadd_bw__read;
  wire [512:0] qr26_vadd_bw__din;
  wire qr26_vadd_bw__full_n;
  wire qr26_vadd_bw__write;
  wire [512:0] qr27_vadd_bw__dout;
  wire qr27_vadd_bw__empty_n;
  wire qr27_vadd_bw__read;
  wire [512:0] qr27_vadd_bw__din;
  wire qr27_vadd_bw__full_n;
  wire qr27_vadd_bw__write;
  wire [512:0] qr2_vadd_bw__dout;
  wire qr2_vadd_bw__empty_n;
  wire qr2_vadd_bw__read;
  wire [512:0] qr2_vadd_bw__din;
  wire qr2_vadd_bw__full_n;
  wire qr2_vadd_bw__write;
  wire [512:0] qr3_vadd_bw__dout;
  wire qr3_vadd_bw__empty_n;
  wire qr3_vadd_bw__read;
  wire [512:0] qr3_vadd_bw__din;
  wire qr3_vadd_bw__full_n;
  wire qr3_vadd_bw__write;
  wire [512:0] qr4_vadd_bw__dout;
  wire qr4_vadd_bw__empty_n;
  wire qr4_vadd_bw__read;
  wire [512:0] qr4_vadd_bw__din;
  wire qr4_vadd_bw__full_n;
  wire qr4_vadd_bw__write;
  wire [512:0] qr5_vadd_bw__dout;
  wire qr5_vadd_bw__empty_n;
  wire qr5_vadd_bw__read;
  wire [512:0] qr5_vadd_bw__din;
  wire qr5_vadd_bw__full_n;
  wire qr5_vadd_bw__write;
  wire [512:0] qr6_vadd_bw__dout;
  wire qr6_vadd_bw__empty_n;
  wire qr6_vadd_bw__read;
  wire [512:0] qr6_vadd_bw__din;
  wire qr6_vadd_bw__full_n;
  wire qr6_vadd_bw__write;
  wire [512:0] qr7_vadd_bw__dout;
  wire qr7_vadd_bw__empty_n;
  wire qr7_vadd_bw__read;
  wire [512:0] qr7_vadd_bw__din;
  wire qr7_vadd_bw__full_n;
  wire qr7_vadd_bw__write;
  wire [512:0] qr8_vadd_bw__dout;
  wire qr8_vadd_bw__empty_n;
  wire qr8_vadd_bw__read;
  wire [512:0] qr8_vadd_bw__din;
  wire qr8_vadd_bw__full_n;
  wire qr8_vadd_bw__write;
  wire [512:0] qr9_vadd_bw__dout;
  wire qr9_vadd_bw__empty_n;
  wire qr9_vadd_bw__read;
  wire [512:0] qr9_vadd_bw__din;
  wire qr9_vadd_bw__full_n;
  wire qr9_vadd_bw__write;
  wire [512:0] qw0_vadd_bw__dout;
  wire qw0_vadd_bw__empty_n;
  wire qw0_vadd_bw__read;
  wire [512:0] qw0_vadd_bw__din;
  wire qw0_vadd_bw__full_n;
  wire qw0_vadd_bw__write;
  wire [512:0] qw10_vadd_bw__dout;
  wire qw10_vadd_bw__empty_n;
  wire qw10_vadd_bw__read;
  wire [512:0] qw10_vadd_bw__din;
  wire qw10_vadd_bw__full_n;
  wire qw10_vadd_bw__write;
  wire [512:0] qw11_vadd_bw__dout;
  wire qw11_vadd_bw__empty_n;
  wire qw11_vadd_bw__read;
  wire [512:0] qw11_vadd_bw__din;
  wire qw11_vadd_bw__full_n;
  wire qw11_vadd_bw__write;
  wire [512:0] qw12_vadd_bw__dout;
  wire qw12_vadd_bw__empty_n;
  wire qw12_vadd_bw__read;
  wire [512:0] qw12_vadd_bw__din;
  wire qw12_vadd_bw__full_n;
  wire qw12_vadd_bw__write;
  wire [512:0] qw13_vadd_bw__dout;
  wire qw13_vadd_bw__empty_n;
  wire qw13_vadd_bw__read;
  wire [512:0] qw13_vadd_bw__din;
  wire qw13_vadd_bw__full_n;
  wire qw13_vadd_bw__write;
  wire [512:0] qw14_vadd_bw__dout;
  wire qw14_vadd_bw__empty_n;
  wire qw14_vadd_bw__read;
  wire [512:0] qw14_vadd_bw__din;
  wire qw14_vadd_bw__full_n;
  wire qw14_vadd_bw__write;
  wire [512:0] qw15_vadd_bw__dout;
  wire qw15_vadd_bw__empty_n;
  wire qw15_vadd_bw__read;
  wire [512:0] qw15_vadd_bw__din;
  wire qw15_vadd_bw__full_n;
  wire qw15_vadd_bw__write;
  wire [512:0] qw16_vadd_bw__dout;
  wire qw16_vadd_bw__empty_n;
  wire qw16_vadd_bw__read;
  wire [512:0] qw16_vadd_bw__din;
  wire qw16_vadd_bw__full_n;
  wire qw16_vadd_bw__write;
  wire [512:0] qw17_vadd_bw__dout;
  wire qw17_vadd_bw__empty_n;
  wire qw17_vadd_bw__read;
  wire [512:0] qw17_vadd_bw__din;
  wire qw17_vadd_bw__full_n;
  wire qw17_vadd_bw__write;
  wire [512:0] qw18_vadd_bw__dout;
  wire qw18_vadd_bw__empty_n;
  wire qw18_vadd_bw__read;
  wire [512:0] qw18_vadd_bw__din;
  wire qw18_vadd_bw__full_n;
  wire qw18_vadd_bw__write;
  wire [512:0] qw19_vadd_bw__dout;
  wire qw19_vadd_bw__empty_n;
  wire qw19_vadd_bw__read;
  wire [512:0] qw19_vadd_bw__din;
  wire qw19_vadd_bw__full_n;
  wire qw19_vadd_bw__write;
  wire [512:0] qw1_vadd_bw__dout;
  wire qw1_vadd_bw__empty_n;
  wire qw1_vadd_bw__read;
  wire [512:0] qw1_vadd_bw__din;
  wire qw1_vadd_bw__full_n;
  wire qw1_vadd_bw__write;
  wire [512:0] qw20_vadd_bw__dout;
  wire qw20_vadd_bw__empty_n;
  wire qw20_vadd_bw__read;
  wire [512:0] qw20_vadd_bw__din;
  wire qw20_vadd_bw__full_n;
  wire qw20_vadd_bw__write;
  wire [512:0] qw21_vadd_bw__dout;
  wire qw21_vadd_bw__empty_n;
  wire qw21_vadd_bw__read;
  wire [512:0] qw21_vadd_bw__din;
  wire qw21_vadd_bw__full_n;
  wire qw21_vadd_bw__write;
  wire [512:0] qw22_vadd_bw__dout;
  wire qw22_vadd_bw__empty_n;
  wire qw22_vadd_bw__read;
  wire [512:0] qw22_vadd_bw__din;
  wire qw22_vadd_bw__full_n;
  wire qw22_vadd_bw__write;
  wire [512:0] qw23_vadd_bw__dout;
  wire qw23_vadd_bw__empty_n;
  wire qw23_vadd_bw__read;
  wire [512:0] qw23_vadd_bw__din;
  wire qw23_vadd_bw__full_n;
  wire qw23_vadd_bw__write;
  wire [512:0] qw24_vadd_bw__dout;
  wire qw24_vadd_bw__empty_n;
  wire qw24_vadd_bw__read;
  wire [512:0] qw24_vadd_bw__din;
  wire qw24_vadd_bw__full_n;
  wire qw24_vadd_bw__write;
  wire [512:0] qw25_vadd_bw__dout;
  wire qw25_vadd_bw__empty_n;
  wire qw25_vadd_bw__read;
  wire [512:0] qw25_vadd_bw__din;
  wire qw25_vadd_bw__full_n;
  wire qw25_vadd_bw__write;
  wire [512:0] qw26_vadd_bw__dout;
  wire qw26_vadd_bw__empty_n;
  wire qw26_vadd_bw__read;
  wire [512:0] qw26_vadd_bw__din;
  wire qw26_vadd_bw__full_n;
  wire qw26_vadd_bw__write;
  wire [512:0] qw27_vadd_bw__dout;
  wire qw27_vadd_bw__empty_n;
  wire qw27_vadd_bw__read;
  wire [512:0] qw27_vadd_bw__din;
  wire qw27_vadd_bw__full_n;
  wire qw27_vadd_bw__write;
  wire [512:0] qw2_vadd_bw__dout;
  wire qw2_vadd_bw__empty_n;
  wire qw2_vadd_bw__read;
  wire [512:0] qw2_vadd_bw__din;
  wire qw2_vadd_bw__full_n;
  wire qw2_vadd_bw__write;
  wire [512:0] qw3_vadd_bw__dout;
  wire qw3_vadd_bw__empty_n;
  wire qw3_vadd_bw__read;
  wire [512:0] qw3_vadd_bw__din;
  wire qw3_vadd_bw__full_n;
  wire qw3_vadd_bw__write;
  wire [512:0] qw4_vadd_bw__dout;
  wire qw4_vadd_bw__empty_n;
  wire qw4_vadd_bw__read;
  wire [512:0] qw4_vadd_bw__din;
  wire qw4_vadd_bw__full_n;
  wire qw4_vadd_bw__write;
  wire [512:0] qw5_vadd_bw__dout;
  wire qw5_vadd_bw__empty_n;
  wire qw5_vadd_bw__read;
  wire [512:0] qw5_vadd_bw__din;
  wire qw5_vadd_bw__full_n;
  wire qw5_vadd_bw__write;
  wire [512:0] qw6_vadd_bw__dout;
  wire qw6_vadd_bw__empty_n;
  wire qw6_vadd_bw__read;
  wire [512:0] qw6_vadd_bw__din;
  wire qw6_vadd_bw__full_n;
  wire qw6_vadd_bw__write;
  wire [512:0] qw7_vadd_bw__dout;
  wire qw7_vadd_bw__empty_n;
  wire qw7_vadd_bw__read;
  wire [512:0] qw7_vadd_bw__din;
  wire qw7_vadd_bw__full_n;
  wire qw7_vadd_bw__write;
  wire [512:0] qw8_vadd_bw__dout;
  wire qw8_vadd_bw__empty_n;
  wire qw8_vadd_bw__read;
  wire [512:0] qw8_vadd_bw__din;
  wire qw8_vadd_bw__full_n;
  wire qw8_vadd_bw__write;
  wire [512:0] qw9_vadd_bw__dout;
  wire qw9_vadd_bw__empty_n;
  wire qw9_vadd_bw__read;
  wire [512:0] qw9_vadd_bw__din;
  wire qw9_vadd_bw__full_n;
  wire qw9_vadd_bw__write;
  wire [63:0] m_axi_rmem0___Mmap2Stream_0___mmap_ARADDR;
  wire [1:0] m_axi_rmem0___Mmap2Stream_0___mmap_ARBURST;
  wire [3:0] m_axi_rmem0___Mmap2Stream_0___mmap_ARCACHE;
  wire [0:0] m_axi_rmem0___Mmap2Stream_0___mmap_ARID;
  wire [7:0] m_axi_rmem0___Mmap2Stream_0___mmap_ARLEN;
  wire m_axi_rmem0___Mmap2Stream_0___mmap_ARLOCK;
  wire [2:0] m_axi_rmem0___Mmap2Stream_0___mmap_ARPROT;
  wire [3:0] m_axi_rmem0___Mmap2Stream_0___mmap_ARQOS;
  wire m_axi_rmem0___Mmap2Stream_0___mmap_ARREADY;
  wire [2:0] m_axi_rmem0___Mmap2Stream_0___mmap_ARSIZE;
  wire m_axi_rmem0___Mmap2Stream_0___mmap_ARVALID;
  wire [63:0] m_axi_rmem0___Mmap2Stream_0___mmap_AWADDR;
  wire [1:0] m_axi_rmem0___Mmap2Stream_0___mmap_AWBURST;
  wire [3:0] m_axi_rmem0___Mmap2Stream_0___mmap_AWCACHE;
  wire [0:0] m_axi_rmem0___Mmap2Stream_0___mmap_AWID;
  wire [7:0] m_axi_rmem0___Mmap2Stream_0___mmap_AWLEN;
  wire m_axi_rmem0___Mmap2Stream_0___mmap_AWLOCK;
  wire [2:0] m_axi_rmem0___Mmap2Stream_0___mmap_AWPROT;
  wire [3:0] m_axi_rmem0___Mmap2Stream_0___mmap_AWQOS;
  wire m_axi_rmem0___Mmap2Stream_0___mmap_AWREADY;
  wire [2:0] m_axi_rmem0___Mmap2Stream_0___mmap_AWSIZE;
  wire m_axi_rmem0___Mmap2Stream_0___mmap_AWVALID;
  wire [0:0] m_axi_rmem0___Mmap2Stream_0___mmap_BID;
  wire m_axi_rmem0___Mmap2Stream_0___mmap_BREADY;
  wire [1:0] m_axi_rmem0___Mmap2Stream_0___mmap_BRESP;
  wire m_axi_rmem0___Mmap2Stream_0___mmap_BVALID;
  wire [511:0] m_axi_rmem0___Mmap2Stream_0___mmap_RDATA;
  wire [0:0] m_axi_rmem0___Mmap2Stream_0___mmap_RID;
  wire m_axi_rmem0___Mmap2Stream_0___mmap_RLAST;
  wire m_axi_rmem0___Mmap2Stream_0___mmap_RREADY;
  wire [1:0] m_axi_rmem0___Mmap2Stream_0___mmap_RRESP;
  wire m_axi_rmem0___Mmap2Stream_0___mmap_RVALID;
  wire [511:0] m_axi_rmem0___Mmap2Stream_0___mmap_WDATA;
  wire m_axi_rmem0___Mmap2Stream_0___mmap_WLAST;
  wire m_axi_rmem0___Mmap2Stream_0___mmap_WREADY;
  wire [63:0] m_axi_rmem0___Mmap2Stream_0___mmap_WSTRB;
  wire m_axi_rmem0___Mmap2Stream_0___mmap_WVALID;
  wire [63:0] m_axi_rmem0___Stream2Mmap_0___mmap_ARADDR;
  wire [1:0] m_axi_rmem0___Stream2Mmap_0___mmap_ARBURST;
  wire [3:0] m_axi_rmem0___Stream2Mmap_0___mmap_ARCACHE;
  wire [0:0] m_axi_rmem0___Stream2Mmap_0___mmap_ARID;
  wire [7:0] m_axi_rmem0___Stream2Mmap_0___mmap_ARLEN;
  wire m_axi_rmem0___Stream2Mmap_0___mmap_ARLOCK;
  wire [2:0] m_axi_rmem0___Stream2Mmap_0___mmap_ARPROT;
  wire [3:0] m_axi_rmem0___Stream2Mmap_0___mmap_ARQOS;
  wire m_axi_rmem0___Stream2Mmap_0___mmap_ARREADY;
  wire [2:0] m_axi_rmem0___Stream2Mmap_0___mmap_ARSIZE;
  wire m_axi_rmem0___Stream2Mmap_0___mmap_ARVALID;
  wire [63:0] m_axi_rmem0___Stream2Mmap_0___mmap_AWADDR;
  wire [1:0] m_axi_rmem0___Stream2Mmap_0___mmap_AWBURST;
  wire [3:0] m_axi_rmem0___Stream2Mmap_0___mmap_AWCACHE;
  wire [0:0] m_axi_rmem0___Stream2Mmap_0___mmap_AWID;
  wire [7:0] m_axi_rmem0___Stream2Mmap_0___mmap_AWLEN;
  wire m_axi_rmem0___Stream2Mmap_0___mmap_AWLOCK;
  wire [2:0] m_axi_rmem0___Stream2Mmap_0___mmap_AWPROT;
  wire [3:0] m_axi_rmem0___Stream2Mmap_0___mmap_AWQOS;
  wire m_axi_rmem0___Stream2Mmap_0___mmap_AWREADY;
  wire [2:0] m_axi_rmem0___Stream2Mmap_0___mmap_AWSIZE;
  wire m_axi_rmem0___Stream2Mmap_0___mmap_AWVALID;
  wire [0:0] m_axi_rmem0___Stream2Mmap_0___mmap_BID;
  wire m_axi_rmem0___Stream2Mmap_0___mmap_BREADY;
  wire [1:0] m_axi_rmem0___Stream2Mmap_0___mmap_BRESP;
  wire m_axi_rmem0___Stream2Mmap_0___mmap_BVALID;
  wire [511:0] m_axi_rmem0___Stream2Mmap_0___mmap_RDATA;
  wire [0:0] m_axi_rmem0___Stream2Mmap_0___mmap_RID;
  wire m_axi_rmem0___Stream2Mmap_0___mmap_RLAST;
  wire m_axi_rmem0___Stream2Mmap_0___mmap_RREADY;
  wire [1:0] m_axi_rmem0___Stream2Mmap_0___mmap_RRESP;
  wire m_axi_rmem0___Stream2Mmap_0___mmap_RVALID;
  wire [511:0] m_axi_rmem0___Stream2Mmap_0___mmap_WDATA;
  wire m_axi_rmem0___Stream2Mmap_0___mmap_WLAST;
  wire m_axi_rmem0___Stream2Mmap_0___mmap_WREADY;
  wire [63:0] m_axi_rmem0___Stream2Mmap_0___mmap_WSTRB;
  wire m_axi_rmem0___Stream2Mmap_0___mmap_WVALID;
  wire [63:0] m_axi_rmem1___Mmap2Stream_1___mmap_ARADDR;
  wire [1:0] m_axi_rmem1___Mmap2Stream_1___mmap_ARBURST;
  wire [3:0] m_axi_rmem1___Mmap2Stream_1___mmap_ARCACHE;
  wire [0:0] m_axi_rmem1___Mmap2Stream_1___mmap_ARID;
  wire [7:0] m_axi_rmem1___Mmap2Stream_1___mmap_ARLEN;
  wire m_axi_rmem1___Mmap2Stream_1___mmap_ARLOCK;
  wire [2:0] m_axi_rmem1___Mmap2Stream_1___mmap_ARPROT;
  wire [3:0] m_axi_rmem1___Mmap2Stream_1___mmap_ARQOS;
  wire m_axi_rmem1___Mmap2Stream_1___mmap_ARREADY;
  wire [2:0] m_axi_rmem1___Mmap2Stream_1___mmap_ARSIZE;
  wire m_axi_rmem1___Mmap2Stream_1___mmap_ARVALID;
  wire [63:0] m_axi_rmem1___Mmap2Stream_1___mmap_AWADDR;
  wire [1:0] m_axi_rmem1___Mmap2Stream_1___mmap_AWBURST;
  wire [3:0] m_axi_rmem1___Mmap2Stream_1___mmap_AWCACHE;
  wire [0:0] m_axi_rmem1___Mmap2Stream_1___mmap_AWID;
  wire [7:0] m_axi_rmem1___Mmap2Stream_1___mmap_AWLEN;
  wire m_axi_rmem1___Mmap2Stream_1___mmap_AWLOCK;
  wire [2:0] m_axi_rmem1___Mmap2Stream_1___mmap_AWPROT;
  wire [3:0] m_axi_rmem1___Mmap2Stream_1___mmap_AWQOS;
  wire m_axi_rmem1___Mmap2Stream_1___mmap_AWREADY;
  wire [2:0] m_axi_rmem1___Mmap2Stream_1___mmap_AWSIZE;
  wire m_axi_rmem1___Mmap2Stream_1___mmap_AWVALID;
  wire [0:0] m_axi_rmem1___Mmap2Stream_1___mmap_BID;
  wire m_axi_rmem1___Mmap2Stream_1___mmap_BREADY;
  wire [1:0] m_axi_rmem1___Mmap2Stream_1___mmap_BRESP;
  wire m_axi_rmem1___Mmap2Stream_1___mmap_BVALID;
  wire [511:0] m_axi_rmem1___Mmap2Stream_1___mmap_RDATA;
  wire [0:0] m_axi_rmem1___Mmap2Stream_1___mmap_RID;
  wire m_axi_rmem1___Mmap2Stream_1___mmap_RLAST;
  wire m_axi_rmem1___Mmap2Stream_1___mmap_RREADY;
  wire [1:0] m_axi_rmem1___Mmap2Stream_1___mmap_RRESP;
  wire m_axi_rmem1___Mmap2Stream_1___mmap_RVALID;
  wire [511:0] m_axi_rmem1___Mmap2Stream_1___mmap_WDATA;
  wire m_axi_rmem1___Mmap2Stream_1___mmap_WLAST;
  wire m_axi_rmem1___Mmap2Stream_1___mmap_WREADY;
  wire [63:0] m_axi_rmem1___Mmap2Stream_1___mmap_WSTRB;
  wire m_axi_rmem1___Mmap2Stream_1___mmap_WVALID;
  wire [63:0] m_axi_rmem1___Stream2Mmap_1___mmap_ARADDR;
  wire [1:0] m_axi_rmem1___Stream2Mmap_1___mmap_ARBURST;
  wire [3:0] m_axi_rmem1___Stream2Mmap_1___mmap_ARCACHE;
  wire [0:0] m_axi_rmem1___Stream2Mmap_1___mmap_ARID;
  wire [7:0] m_axi_rmem1___Stream2Mmap_1___mmap_ARLEN;
  wire m_axi_rmem1___Stream2Mmap_1___mmap_ARLOCK;
  wire [2:0] m_axi_rmem1___Stream2Mmap_1___mmap_ARPROT;
  wire [3:0] m_axi_rmem1___Stream2Mmap_1___mmap_ARQOS;
  wire m_axi_rmem1___Stream2Mmap_1___mmap_ARREADY;
  wire [2:0] m_axi_rmem1___Stream2Mmap_1___mmap_ARSIZE;
  wire m_axi_rmem1___Stream2Mmap_1___mmap_ARVALID;
  wire [63:0] m_axi_rmem1___Stream2Mmap_1___mmap_AWADDR;
  wire [1:0] m_axi_rmem1___Stream2Mmap_1___mmap_AWBURST;
  wire [3:0] m_axi_rmem1___Stream2Mmap_1___mmap_AWCACHE;
  wire [0:0] m_axi_rmem1___Stream2Mmap_1___mmap_AWID;
  wire [7:0] m_axi_rmem1___Stream2Mmap_1___mmap_AWLEN;
  wire m_axi_rmem1___Stream2Mmap_1___mmap_AWLOCK;
  wire [2:0] m_axi_rmem1___Stream2Mmap_1___mmap_AWPROT;
  wire [3:0] m_axi_rmem1___Stream2Mmap_1___mmap_AWQOS;
  wire m_axi_rmem1___Stream2Mmap_1___mmap_AWREADY;
  wire [2:0] m_axi_rmem1___Stream2Mmap_1___mmap_AWSIZE;
  wire m_axi_rmem1___Stream2Mmap_1___mmap_AWVALID;
  wire [0:0] m_axi_rmem1___Stream2Mmap_1___mmap_BID;
  wire m_axi_rmem1___Stream2Mmap_1___mmap_BREADY;
  wire [1:0] m_axi_rmem1___Stream2Mmap_1___mmap_BRESP;
  wire m_axi_rmem1___Stream2Mmap_1___mmap_BVALID;
  wire [511:0] m_axi_rmem1___Stream2Mmap_1___mmap_RDATA;
  wire [0:0] m_axi_rmem1___Stream2Mmap_1___mmap_RID;
  wire m_axi_rmem1___Stream2Mmap_1___mmap_RLAST;
  wire m_axi_rmem1___Stream2Mmap_1___mmap_RREADY;
  wire [1:0] m_axi_rmem1___Stream2Mmap_1___mmap_RRESP;
  wire m_axi_rmem1___Stream2Mmap_1___mmap_RVALID;
  wire [511:0] m_axi_rmem1___Stream2Mmap_1___mmap_WDATA;
  wire m_axi_rmem1___Stream2Mmap_1___mmap_WLAST;
  wire m_axi_rmem1___Stream2Mmap_1___mmap_WREADY;
  wire [63:0] m_axi_rmem1___Stream2Mmap_1___mmap_WSTRB;
  wire m_axi_rmem1___Stream2Mmap_1___mmap_WVALID;
  wire [63:0] m_axi_rmem2___Mmap2Stream_2___mmap_ARADDR;
  wire [1:0] m_axi_rmem2___Mmap2Stream_2___mmap_ARBURST;
  wire [3:0] m_axi_rmem2___Mmap2Stream_2___mmap_ARCACHE;
  wire [0:0] m_axi_rmem2___Mmap2Stream_2___mmap_ARID;
  wire [7:0] m_axi_rmem2___Mmap2Stream_2___mmap_ARLEN;
  wire m_axi_rmem2___Mmap2Stream_2___mmap_ARLOCK;
  wire [2:0] m_axi_rmem2___Mmap2Stream_2___mmap_ARPROT;
  wire [3:0] m_axi_rmem2___Mmap2Stream_2___mmap_ARQOS;
  wire m_axi_rmem2___Mmap2Stream_2___mmap_ARREADY;
  wire [2:0] m_axi_rmem2___Mmap2Stream_2___mmap_ARSIZE;
  wire m_axi_rmem2___Mmap2Stream_2___mmap_ARVALID;
  wire [63:0] m_axi_rmem2___Mmap2Stream_2___mmap_AWADDR;
  wire [1:0] m_axi_rmem2___Mmap2Stream_2___mmap_AWBURST;
  wire [3:0] m_axi_rmem2___Mmap2Stream_2___mmap_AWCACHE;
  wire [0:0] m_axi_rmem2___Mmap2Stream_2___mmap_AWID;
  wire [7:0] m_axi_rmem2___Mmap2Stream_2___mmap_AWLEN;
  wire m_axi_rmem2___Mmap2Stream_2___mmap_AWLOCK;
  wire [2:0] m_axi_rmem2___Mmap2Stream_2___mmap_AWPROT;
  wire [3:0] m_axi_rmem2___Mmap2Stream_2___mmap_AWQOS;
  wire m_axi_rmem2___Mmap2Stream_2___mmap_AWREADY;
  wire [2:0] m_axi_rmem2___Mmap2Stream_2___mmap_AWSIZE;
  wire m_axi_rmem2___Mmap2Stream_2___mmap_AWVALID;
  wire [0:0] m_axi_rmem2___Mmap2Stream_2___mmap_BID;
  wire m_axi_rmem2___Mmap2Stream_2___mmap_BREADY;
  wire [1:0] m_axi_rmem2___Mmap2Stream_2___mmap_BRESP;
  wire m_axi_rmem2___Mmap2Stream_2___mmap_BVALID;
  wire [511:0] m_axi_rmem2___Mmap2Stream_2___mmap_RDATA;
  wire [0:0] m_axi_rmem2___Mmap2Stream_2___mmap_RID;
  wire m_axi_rmem2___Mmap2Stream_2___mmap_RLAST;
  wire m_axi_rmem2___Mmap2Stream_2___mmap_RREADY;
  wire [1:0] m_axi_rmem2___Mmap2Stream_2___mmap_RRESP;
  wire m_axi_rmem2___Mmap2Stream_2___mmap_RVALID;
  wire [511:0] m_axi_rmem2___Mmap2Stream_2___mmap_WDATA;
  wire m_axi_rmem2___Mmap2Stream_2___mmap_WLAST;
  wire m_axi_rmem2___Mmap2Stream_2___mmap_WREADY;
  wire [63:0] m_axi_rmem2___Mmap2Stream_2___mmap_WSTRB;
  wire m_axi_rmem2___Mmap2Stream_2___mmap_WVALID;
  wire [63:0] m_axi_rmem2___Stream2Mmap_2___mmap_ARADDR;
  wire [1:0] m_axi_rmem2___Stream2Mmap_2___mmap_ARBURST;
  wire [3:0] m_axi_rmem2___Stream2Mmap_2___mmap_ARCACHE;
  wire [0:0] m_axi_rmem2___Stream2Mmap_2___mmap_ARID;
  wire [7:0] m_axi_rmem2___Stream2Mmap_2___mmap_ARLEN;
  wire m_axi_rmem2___Stream2Mmap_2___mmap_ARLOCK;
  wire [2:0] m_axi_rmem2___Stream2Mmap_2___mmap_ARPROT;
  wire [3:0] m_axi_rmem2___Stream2Mmap_2___mmap_ARQOS;
  wire m_axi_rmem2___Stream2Mmap_2___mmap_ARREADY;
  wire [2:0] m_axi_rmem2___Stream2Mmap_2___mmap_ARSIZE;
  wire m_axi_rmem2___Stream2Mmap_2___mmap_ARVALID;
  wire [63:0] m_axi_rmem2___Stream2Mmap_2___mmap_AWADDR;
  wire [1:0] m_axi_rmem2___Stream2Mmap_2___mmap_AWBURST;
  wire [3:0] m_axi_rmem2___Stream2Mmap_2___mmap_AWCACHE;
  wire [0:0] m_axi_rmem2___Stream2Mmap_2___mmap_AWID;
  wire [7:0] m_axi_rmem2___Stream2Mmap_2___mmap_AWLEN;
  wire m_axi_rmem2___Stream2Mmap_2___mmap_AWLOCK;
  wire [2:0] m_axi_rmem2___Stream2Mmap_2___mmap_AWPROT;
  wire [3:0] m_axi_rmem2___Stream2Mmap_2___mmap_AWQOS;
  wire m_axi_rmem2___Stream2Mmap_2___mmap_AWREADY;
  wire [2:0] m_axi_rmem2___Stream2Mmap_2___mmap_AWSIZE;
  wire m_axi_rmem2___Stream2Mmap_2___mmap_AWVALID;
  wire [0:0] m_axi_rmem2___Stream2Mmap_2___mmap_BID;
  wire m_axi_rmem2___Stream2Mmap_2___mmap_BREADY;
  wire [1:0] m_axi_rmem2___Stream2Mmap_2___mmap_BRESP;
  wire m_axi_rmem2___Stream2Mmap_2___mmap_BVALID;
  wire [511:0] m_axi_rmem2___Stream2Mmap_2___mmap_RDATA;
  wire [0:0] m_axi_rmem2___Stream2Mmap_2___mmap_RID;
  wire m_axi_rmem2___Stream2Mmap_2___mmap_RLAST;
  wire m_axi_rmem2___Stream2Mmap_2___mmap_RREADY;
  wire [1:0] m_axi_rmem2___Stream2Mmap_2___mmap_RRESP;
  wire m_axi_rmem2___Stream2Mmap_2___mmap_RVALID;
  wire [511:0] m_axi_rmem2___Stream2Mmap_2___mmap_WDATA;
  wire m_axi_rmem2___Stream2Mmap_2___mmap_WLAST;
  wire m_axi_rmem2___Stream2Mmap_2___mmap_WREADY;
  wire [63:0] m_axi_rmem2___Stream2Mmap_2___mmap_WSTRB;
  wire m_axi_rmem2___Stream2Mmap_2___mmap_WVALID;
  wire [63:0] m_axi_rmem3___Mmap2Stream_3___mmap_ARADDR;
  wire [1:0] m_axi_rmem3___Mmap2Stream_3___mmap_ARBURST;
  wire [3:0] m_axi_rmem3___Mmap2Stream_3___mmap_ARCACHE;
  wire [0:0] m_axi_rmem3___Mmap2Stream_3___mmap_ARID;
  wire [7:0] m_axi_rmem3___Mmap2Stream_3___mmap_ARLEN;
  wire m_axi_rmem3___Mmap2Stream_3___mmap_ARLOCK;
  wire [2:0] m_axi_rmem3___Mmap2Stream_3___mmap_ARPROT;
  wire [3:0] m_axi_rmem3___Mmap2Stream_3___mmap_ARQOS;
  wire m_axi_rmem3___Mmap2Stream_3___mmap_ARREADY;
  wire [2:0] m_axi_rmem3___Mmap2Stream_3___mmap_ARSIZE;
  wire m_axi_rmem3___Mmap2Stream_3___mmap_ARVALID;
  wire [63:0] m_axi_rmem3___Mmap2Stream_3___mmap_AWADDR;
  wire [1:0] m_axi_rmem3___Mmap2Stream_3___mmap_AWBURST;
  wire [3:0] m_axi_rmem3___Mmap2Stream_3___mmap_AWCACHE;
  wire [0:0] m_axi_rmem3___Mmap2Stream_3___mmap_AWID;
  wire [7:0] m_axi_rmem3___Mmap2Stream_3___mmap_AWLEN;
  wire m_axi_rmem3___Mmap2Stream_3___mmap_AWLOCK;
  wire [2:0] m_axi_rmem3___Mmap2Stream_3___mmap_AWPROT;
  wire [3:0] m_axi_rmem3___Mmap2Stream_3___mmap_AWQOS;
  wire m_axi_rmem3___Mmap2Stream_3___mmap_AWREADY;
  wire [2:0] m_axi_rmem3___Mmap2Stream_3___mmap_AWSIZE;
  wire m_axi_rmem3___Mmap2Stream_3___mmap_AWVALID;
  wire [0:0] m_axi_rmem3___Mmap2Stream_3___mmap_BID;
  wire m_axi_rmem3___Mmap2Stream_3___mmap_BREADY;
  wire [1:0] m_axi_rmem3___Mmap2Stream_3___mmap_BRESP;
  wire m_axi_rmem3___Mmap2Stream_3___mmap_BVALID;
  wire [511:0] m_axi_rmem3___Mmap2Stream_3___mmap_RDATA;
  wire [0:0] m_axi_rmem3___Mmap2Stream_3___mmap_RID;
  wire m_axi_rmem3___Mmap2Stream_3___mmap_RLAST;
  wire m_axi_rmem3___Mmap2Stream_3___mmap_RREADY;
  wire [1:0] m_axi_rmem3___Mmap2Stream_3___mmap_RRESP;
  wire m_axi_rmem3___Mmap2Stream_3___mmap_RVALID;
  wire [511:0] m_axi_rmem3___Mmap2Stream_3___mmap_WDATA;
  wire m_axi_rmem3___Mmap2Stream_3___mmap_WLAST;
  wire m_axi_rmem3___Mmap2Stream_3___mmap_WREADY;
  wire [63:0] m_axi_rmem3___Mmap2Stream_3___mmap_WSTRB;
  wire m_axi_rmem3___Mmap2Stream_3___mmap_WVALID;
  wire [63:0] m_axi_rmem3___Stream2Mmap_3___mmap_ARADDR;
  wire [1:0] m_axi_rmem3___Stream2Mmap_3___mmap_ARBURST;
  wire [3:0] m_axi_rmem3___Stream2Mmap_3___mmap_ARCACHE;
  wire [0:0] m_axi_rmem3___Stream2Mmap_3___mmap_ARID;
  wire [7:0] m_axi_rmem3___Stream2Mmap_3___mmap_ARLEN;
  wire m_axi_rmem3___Stream2Mmap_3___mmap_ARLOCK;
  wire [2:0] m_axi_rmem3___Stream2Mmap_3___mmap_ARPROT;
  wire [3:0] m_axi_rmem3___Stream2Mmap_3___mmap_ARQOS;
  wire m_axi_rmem3___Stream2Mmap_3___mmap_ARREADY;
  wire [2:0] m_axi_rmem3___Stream2Mmap_3___mmap_ARSIZE;
  wire m_axi_rmem3___Stream2Mmap_3___mmap_ARVALID;
  wire [63:0] m_axi_rmem3___Stream2Mmap_3___mmap_AWADDR;
  wire [1:0] m_axi_rmem3___Stream2Mmap_3___mmap_AWBURST;
  wire [3:0] m_axi_rmem3___Stream2Mmap_3___mmap_AWCACHE;
  wire [0:0] m_axi_rmem3___Stream2Mmap_3___mmap_AWID;
  wire [7:0] m_axi_rmem3___Stream2Mmap_3___mmap_AWLEN;
  wire m_axi_rmem3___Stream2Mmap_3___mmap_AWLOCK;
  wire [2:0] m_axi_rmem3___Stream2Mmap_3___mmap_AWPROT;
  wire [3:0] m_axi_rmem3___Stream2Mmap_3___mmap_AWQOS;
  wire m_axi_rmem3___Stream2Mmap_3___mmap_AWREADY;
  wire [2:0] m_axi_rmem3___Stream2Mmap_3___mmap_AWSIZE;
  wire m_axi_rmem3___Stream2Mmap_3___mmap_AWVALID;
  wire [0:0] m_axi_rmem3___Stream2Mmap_3___mmap_BID;
  wire m_axi_rmem3___Stream2Mmap_3___mmap_BREADY;
  wire [1:0] m_axi_rmem3___Stream2Mmap_3___mmap_BRESP;
  wire m_axi_rmem3___Stream2Mmap_3___mmap_BVALID;
  wire [511:0] m_axi_rmem3___Stream2Mmap_3___mmap_RDATA;
  wire [0:0] m_axi_rmem3___Stream2Mmap_3___mmap_RID;
  wire m_axi_rmem3___Stream2Mmap_3___mmap_RLAST;
  wire m_axi_rmem3___Stream2Mmap_3___mmap_RREADY;
  wire [1:0] m_axi_rmem3___Stream2Mmap_3___mmap_RRESP;
  wire m_axi_rmem3___Stream2Mmap_3___mmap_RVALID;
  wire [511:0] m_axi_rmem3___Stream2Mmap_3___mmap_WDATA;
  wire m_axi_rmem3___Stream2Mmap_3___mmap_WLAST;
  wire m_axi_rmem3___Stream2Mmap_3___mmap_WREADY;
  wire [63:0] m_axi_rmem3___Stream2Mmap_3___mmap_WSTRB;
  wire m_axi_rmem3___Stream2Mmap_3___mmap_WVALID;
  wire [63:0] m_axi_rmem4___Mmap2Stream_4___mmap_ARADDR;
  wire [1:0] m_axi_rmem4___Mmap2Stream_4___mmap_ARBURST;
  wire [3:0] m_axi_rmem4___Mmap2Stream_4___mmap_ARCACHE;
  wire [0:0] m_axi_rmem4___Mmap2Stream_4___mmap_ARID;
  wire [7:0] m_axi_rmem4___Mmap2Stream_4___mmap_ARLEN;
  wire m_axi_rmem4___Mmap2Stream_4___mmap_ARLOCK;
  wire [2:0] m_axi_rmem4___Mmap2Stream_4___mmap_ARPROT;
  wire [3:0] m_axi_rmem4___Mmap2Stream_4___mmap_ARQOS;
  wire m_axi_rmem4___Mmap2Stream_4___mmap_ARREADY;
  wire [2:0] m_axi_rmem4___Mmap2Stream_4___mmap_ARSIZE;
  wire m_axi_rmem4___Mmap2Stream_4___mmap_ARVALID;
  wire [63:0] m_axi_rmem4___Mmap2Stream_4___mmap_AWADDR;
  wire [1:0] m_axi_rmem4___Mmap2Stream_4___mmap_AWBURST;
  wire [3:0] m_axi_rmem4___Mmap2Stream_4___mmap_AWCACHE;
  wire [0:0] m_axi_rmem4___Mmap2Stream_4___mmap_AWID;
  wire [7:0] m_axi_rmem4___Mmap2Stream_4___mmap_AWLEN;
  wire m_axi_rmem4___Mmap2Stream_4___mmap_AWLOCK;
  wire [2:0] m_axi_rmem4___Mmap2Stream_4___mmap_AWPROT;
  wire [3:0] m_axi_rmem4___Mmap2Stream_4___mmap_AWQOS;
  wire m_axi_rmem4___Mmap2Stream_4___mmap_AWREADY;
  wire [2:0] m_axi_rmem4___Mmap2Stream_4___mmap_AWSIZE;
  wire m_axi_rmem4___Mmap2Stream_4___mmap_AWVALID;
  wire [0:0] m_axi_rmem4___Mmap2Stream_4___mmap_BID;
  wire m_axi_rmem4___Mmap2Stream_4___mmap_BREADY;
  wire [1:0] m_axi_rmem4___Mmap2Stream_4___mmap_BRESP;
  wire m_axi_rmem4___Mmap2Stream_4___mmap_BVALID;
  wire [511:0] m_axi_rmem4___Mmap2Stream_4___mmap_RDATA;
  wire [0:0] m_axi_rmem4___Mmap2Stream_4___mmap_RID;
  wire m_axi_rmem4___Mmap2Stream_4___mmap_RLAST;
  wire m_axi_rmem4___Mmap2Stream_4___mmap_RREADY;
  wire [1:0] m_axi_rmem4___Mmap2Stream_4___mmap_RRESP;
  wire m_axi_rmem4___Mmap2Stream_4___mmap_RVALID;
  wire [511:0] m_axi_rmem4___Mmap2Stream_4___mmap_WDATA;
  wire m_axi_rmem4___Mmap2Stream_4___mmap_WLAST;
  wire m_axi_rmem4___Mmap2Stream_4___mmap_WREADY;
  wire [63:0] m_axi_rmem4___Mmap2Stream_4___mmap_WSTRB;
  wire m_axi_rmem4___Mmap2Stream_4___mmap_WVALID;
  wire [63:0] m_axi_rmem4___Stream2Mmap_4___mmap_ARADDR;
  wire [1:0] m_axi_rmem4___Stream2Mmap_4___mmap_ARBURST;
  wire [3:0] m_axi_rmem4___Stream2Mmap_4___mmap_ARCACHE;
  wire [0:0] m_axi_rmem4___Stream2Mmap_4___mmap_ARID;
  wire [7:0] m_axi_rmem4___Stream2Mmap_4___mmap_ARLEN;
  wire m_axi_rmem4___Stream2Mmap_4___mmap_ARLOCK;
  wire [2:0] m_axi_rmem4___Stream2Mmap_4___mmap_ARPROT;
  wire [3:0] m_axi_rmem4___Stream2Mmap_4___mmap_ARQOS;
  wire m_axi_rmem4___Stream2Mmap_4___mmap_ARREADY;
  wire [2:0] m_axi_rmem4___Stream2Mmap_4___mmap_ARSIZE;
  wire m_axi_rmem4___Stream2Mmap_4___mmap_ARVALID;
  wire [63:0] m_axi_rmem4___Stream2Mmap_4___mmap_AWADDR;
  wire [1:0] m_axi_rmem4___Stream2Mmap_4___mmap_AWBURST;
  wire [3:0] m_axi_rmem4___Stream2Mmap_4___mmap_AWCACHE;
  wire [0:0] m_axi_rmem4___Stream2Mmap_4___mmap_AWID;
  wire [7:0] m_axi_rmem4___Stream2Mmap_4___mmap_AWLEN;
  wire m_axi_rmem4___Stream2Mmap_4___mmap_AWLOCK;
  wire [2:0] m_axi_rmem4___Stream2Mmap_4___mmap_AWPROT;
  wire [3:0] m_axi_rmem4___Stream2Mmap_4___mmap_AWQOS;
  wire m_axi_rmem4___Stream2Mmap_4___mmap_AWREADY;
  wire [2:0] m_axi_rmem4___Stream2Mmap_4___mmap_AWSIZE;
  wire m_axi_rmem4___Stream2Mmap_4___mmap_AWVALID;
  wire [0:0] m_axi_rmem4___Stream2Mmap_4___mmap_BID;
  wire m_axi_rmem4___Stream2Mmap_4___mmap_BREADY;
  wire [1:0] m_axi_rmem4___Stream2Mmap_4___mmap_BRESP;
  wire m_axi_rmem4___Stream2Mmap_4___mmap_BVALID;
  wire [511:0] m_axi_rmem4___Stream2Mmap_4___mmap_RDATA;
  wire [0:0] m_axi_rmem4___Stream2Mmap_4___mmap_RID;
  wire m_axi_rmem4___Stream2Mmap_4___mmap_RLAST;
  wire m_axi_rmem4___Stream2Mmap_4___mmap_RREADY;
  wire [1:0] m_axi_rmem4___Stream2Mmap_4___mmap_RRESP;
  wire m_axi_rmem4___Stream2Mmap_4___mmap_RVALID;
  wire [511:0] m_axi_rmem4___Stream2Mmap_4___mmap_WDATA;
  wire m_axi_rmem4___Stream2Mmap_4___mmap_WLAST;
  wire m_axi_rmem4___Stream2Mmap_4___mmap_WREADY;
  wire [63:0] m_axi_rmem4___Stream2Mmap_4___mmap_WSTRB;
  wire m_axi_rmem4___Stream2Mmap_4___mmap_WVALID;
  wire [63:0] m_axi_rmem5___Mmap2Stream_5___mmap_ARADDR;
  wire [1:0] m_axi_rmem5___Mmap2Stream_5___mmap_ARBURST;
  wire [3:0] m_axi_rmem5___Mmap2Stream_5___mmap_ARCACHE;
  wire [0:0] m_axi_rmem5___Mmap2Stream_5___mmap_ARID;
  wire [7:0] m_axi_rmem5___Mmap2Stream_5___mmap_ARLEN;
  wire m_axi_rmem5___Mmap2Stream_5___mmap_ARLOCK;
  wire [2:0] m_axi_rmem5___Mmap2Stream_5___mmap_ARPROT;
  wire [3:0] m_axi_rmem5___Mmap2Stream_5___mmap_ARQOS;
  wire m_axi_rmem5___Mmap2Stream_5___mmap_ARREADY;
  wire [2:0] m_axi_rmem5___Mmap2Stream_5___mmap_ARSIZE;
  wire m_axi_rmem5___Mmap2Stream_5___mmap_ARVALID;
  wire [63:0] m_axi_rmem5___Mmap2Stream_5___mmap_AWADDR;
  wire [1:0] m_axi_rmem5___Mmap2Stream_5___mmap_AWBURST;
  wire [3:0] m_axi_rmem5___Mmap2Stream_5___mmap_AWCACHE;
  wire [0:0] m_axi_rmem5___Mmap2Stream_5___mmap_AWID;
  wire [7:0] m_axi_rmem5___Mmap2Stream_5___mmap_AWLEN;
  wire m_axi_rmem5___Mmap2Stream_5___mmap_AWLOCK;
  wire [2:0] m_axi_rmem5___Mmap2Stream_5___mmap_AWPROT;
  wire [3:0] m_axi_rmem5___Mmap2Stream_5___mmap_AWQOS;
  wire m_axi_rmem5___Mmap2Stream_5___mmap_AWREADY;
  wire [2:0] m_axi_rmem5___Mmap2Stream_5___mmap_AWSIZE;
  wire m_axi_rmem5___Mmap2Stream_5___mmap_AWVALID;
  wire [0:0] m_axi_rmem5___Mmap2Stream_5___mmap_BID;
  wire m_axi_rmem5___Mmap2Stream_5___mmap_BREADY;
  wire [1:0] m_axi_rmem5___Mmap2Stream_5___mmap_BRESP;
  wire m_axi_rmem5___Mmap2Stream_5___mmap_BVALID;
  wire [511:0] m_axi_rmem5___Mmap2Stream_5___mmap_RDATA;
  wire [0:0] m_axi_rmem5___Mmap2Stream_5___mmap_RID;
  wire m_axi_rmem5___Mmap2Stream_5___mmap_RLAST;
  wire m_axi_rmem5___Mmap2Stream_5___mmap_RREADY;
  wire [1:0] m_axi_rmem5___Mmap2Stream_5___mmap_RRESP;
  wire m_axi_rmem5___Mmap2Stream_5___mmap_RVALID;
  wire [511:0] m_axi_rmem5___Mmap2Stream_5___mmap_WDATA;
  wire m_axi_rmem5___Mmap2Stream_5___mmap_WLAST;
  wire m_axi_rmem5___Mmap2Stream_5___mmap_WREADY;
  wire [63:0] m_axi_rmem5___Mmap2Stream_5___mmap_WSTRB;
  wire m_axi_rmem5___Mmap2Stream_5___mmap_WVALID;
  wire [63:0] m_axi_rmem5___Stream2Mmap_5___mmap_ARADDR;
  wire [1:0] m_axi_rmem5___Stream2Mmap_5___mmap_ARBURST;
  wire [3:0] m_axi_rmem5___Stream2Mmap_5___mmap_ARCACHE;
  wire [0:0] m_axi_rmem5___Stream2Mmap_5___mmap_ARID;
  wire [7:0] m_axi_rmem5___Stream2Mmap_5___mmap_ARLEN;
  wire m_axi_rmem5___Stream2Mmap_5___mmap_ARLOCK;
  wire [2:0] m_axi_rmem5___Stream2Mmap_5___mmap_ARPROT;
  wire [3:0] m_axi_rmem5___Stream2Mmap_5___mmap_ARQOS;
  wire m_axi_rmem5___Stream2Mmap_5___mmap_ARREADY;
  wire [2:0] m_axi_rmem5___Stream2Mmap_5___mmap_ARSIZE;
  wire m_axi_rmem5___Stream2Mmap_5___mmap_ARVALID;
  wire [63:0] m_axi_rmem5___Stream2Mmap_5___mmap_AWADDR;
  wire [1:0] m_axi_rmem5___Stream2Mmap_5___mmap_AWBURST;
  wire [3:0] m_axi_rmem5___Stream2Mmap_5___mmap_AWCACHE;
  wire [0:0] m_axi_rmem5___Stream2Mmap_5___mmap_AWID;
  wire [7:0] m_axi_rmem5___Stream2Mmap_5___mmap_AWLEN;
  wire m_axi_rmem5___Stream2Mmap_5___mmap_AWLOCK;
  wire [2:0] m_axi_rmem5___Stream2Mmap_5___mmap_AWPROT;
  wire [3:0] m_axi_rmem5___Stream2Mmap_5___mmap_AWQOS;
  wire m_axi_rmem5___Stream2Mmap_5___mmap_AWREADY;
  wire [2:0] m_axi_rmem5___Stream2Mmap_5___mmap_AWSIZE;
  wire m_axi_rmem5___Stream2Mmap_5___mmap_AWVALID;
  wire [0:0] m_axi_rmem5___Stream2Mmap_5___mmap_BID;
  wire m_axi_rmem5___Stream2Mmap_5___mmap_BREADY;
  wire [1:0] m_axi_rmem5___Stream2Mmap_5___mmap_BRESP;
  wire m_axi_rmem5___Stream2Mmap_5___mmap_BVALID;
  wire [511:0] m_axi_rmem5___Stream2Mmap_5___mmap_RDATA;
  wire [0:0] m_axi_rmem5___Stream2Mmap_5___mmap_RID;
  wire m_axi_rmem5___Stream2Mmap_5___mmap_RLAST;
  wire m_axi_rmem5___Stream2Mmap_5___mmap_RREADY;
  wire [1:0] m_axi_rmem5___Stream2Mmap_5___mmap_RRESP;
  wire m_axi_rmem5___Stream2Mmap_5___mmap_RVALID;
  wire [511:0] m_axi_rmem5___Stream2Mmap_5___mmap_WDATA;
  wire m_axi_rmem5___Stream2Mmap_5___mmap_WLAST;
  wire m_axi_rmem5___Stream2Mmap_5___mmap_WREADY;
  wire [63:0] m_axi_rmem5___Stream2Mmap_5___mmap_WSTRB;
  wire m_axi_rmem5___Stream2Mmap_5___mmap_WVALID;
  wire [63:0] m_axi_rmem6___Mmap2Stream_6___mmap_ARADDR;
  wire [1:0] m_axi_rmem6___Mmap2Stream_6___mmap_ARBURST;
  wire [3:0] m_axi_rmem6___Mmap2Stream_6___mmap_ARCACHE;
  wire [0:0] m_axi_rmem6___Mmap2Stream_6___mmap_ARID;
  wire [7:0] m_axi_rmem6___Mmap2Stream_6___mmap_ARLEN;
  wire m_axi_rmem6___Mmap2Stream_6___mmap_ARLOCK;
  wire [2:0] m_axi_rmem6___Mmap2Stream_6___mmap_ARPROT;
  wire [3:0] m_axi_rmem6___Mmap2Stream_6___mmap_ARQOS;
  wire m_axi_rmem6___Mmap2Stream_6___mmap_ARREADY;
  wire [2:0] m_axi_rmem6___Mmap2Stream_6___mmap_ARSIZE;
  wire m_axi_rmem6___Mmap2Stream_6___mmap_ARVALID;
  wire [63:0] m_axi_rmem6___Mmap2Stream_6___mmap_AWADDR;
  wire [1:0] m_axi_rmem6___Mmap2Stream_6___mmap_AWBURST;
  wire [3:0] m_axi_rmem6___Mmap2Stream_6___mmap_AWCACHE;
  wire [0:0] m_axi_rmem6___Mmap2Stream_6___mmap_AWID;
  wire [7:0] m_axi_rmem6___Mmap2Stream_6___mmap_AWLEN;
  wire m_axi_rmem6___Mmap2Stream_6___mmap_AWLOCK;
  wire [2:0] m_axi_rmem6___Mmap2Stream_6___mmap_AWPROT;
  wire [3:0] m_axi_rmem6___Mmap2Stream_6___mmap_AWQOS;
  wire m_axi_rmem6___Mmap2Stream_6___mmap_AWREADY;
  wire [2:0] m_axi_rmem6___Mmap2Stream_6___mmap_AWSIZE;
  wire m_axi_rmem6___Mmap2Stream_6___mmap_AWVALID;
  wire [0:0] m_axi_rmem6___Mmap2Stream_6___mmap_BID;
  wire m_axi_rmem6___Mmap2Stream_6___mmap_BREADY;
  wire [1:0] m_axi_rmem6___Mmap2Stream_6___mmap_BRESP;
  wire m_axi_rmem6___Mmap2Stream_6___mmap_BVALID;
  wire [511:0] m_axi_rmem6___Mmap2Stream_6___mmap_RDATA;
  wire [0:0] m_axi_rmem6___Mmap2Stream_6___mmap_RID;
  wire m_axi_rmem6___Mmap2Stream_6___mmap_RLAST;
  wire m_axi_rmem6___Mmap2Stream_6___mmap_RREADY;
  wire [1:0] m_axi_rmem6___Mmap2Stream_6___mmap_RRESP;
  wire m_axi_rmem6___Mmap2Stream_6___mmap_RVALID;
  wire [511:0] m_axi_rmem6___Mmap2Stream_6___mmap_WDATA;
  wire m_axi_rmem6___Mmap2Stream_6___mmap_WLAST;
  wire m_axi_rmem6___Mmap2Stream_6___mmap_WREADY;
  wire [63:0] m_axi_rmem6___Mmap2Stream_6___mmap_WSTRB;
  wire m_axi_rmem6___Mmap2Stream_6___mmap_WVALID;
  wire [63:0] m_axi_rmem6___Stream2Mmap_6___mmap_ARADDR;
  wire [1:0] m_axi_rmem6___Stream2Mmap_6___mmap_ARBURST;
  wire [3:0] m_axi_rmem6___Stream2Mmap_6___mmap_ARCACHE;
  wire [0:0] m_axi_rmem6___Stream2Mmap_6___mmap_ARID;
  wire [7:0] m_axi_rmem6___Stream2Mmap_6___mmap_ARLEN;
  wire m_axi_rmem6___Stream2Mmap_6___mmap_ARLOCK;
  wire [2:0] m_axi_rmem6___Stream2Mmap_6___mmap_ARPROT;
  wire [3:0] m_axi_rmem6___Stream2Mmap_6___mmap_ARQOS;
  wire m_axi_rmem6___Stream2Mmap_6___mmap_ARREADY;
  wire [2:0] m_axi_rmem6___Stream2Mmap_6___mmap_ARSIZE;
  wire m_axi_rmem6___Stream2Mmap_6___mmap_ARVALID;
  wire [63:0] m_axi_rmem6___Stream2Mmap_6___mmap_AWADDR;
  wire [1:0] m_axi_rmem6___Stream2Mmap_6___mmap_AWBURST;
  wire [3:0] m_axi_rmem6___Stream2Mmap_6___mmap_AWCACHE;
  wire [0:0] m_axi_rmem6___Stream2Mmap_6___mmap_AWID;
  wire [7:0] m_axi_rmem6___Stream2Mmap_6___mmap_AWLEN;
  wire m_axi_rmem6___Stream2Mmap_6___mmap_AWLOCK;
  wire [2:0] m_axi_rmem6___Stream2Mmap_6___mmap_AWPROT;
  wire [3:0] m_axi_rmem6___Stream2Mmap_6___mmap_AWQOS;
  wire m_axi_rmem6___Stream2Mmap_6___mmap_AWREADY;
  wire [2:0] m_axi_rmem6___Stream2Mmap_6___mmap_AWSIZE;
  wire m_axi_rmem6___Stream2Mmap_6___mmap_AWVALID;
  wire [0:0] m_axi_rmem6___Stream2Mmap_6___mmap_BID;
  wire m_axi_rmem6___Stream2Mmap_6___mmap_BREADY;
  wire [1:0] m_axi_rmem6___Stream2Mmap_6___mmap_BRESP;
  wire m_axi_rmem6___Stream2Mmap_6___mmap_BVALID;
  wire [511:0] m_axi_rmem6___Stream2Mmap_6___mmap_RDATA;
  wire [0:0] m_axi_rmem6___Stream2Mmap_6___mmap_RID;
  wire m_axi_rmem6___Stream2Mmap_6___mmap_RLAST;
  wire m_axi_rmem6___Stream2Mmap_6___mmap_RREADY;
  wire [1:0] m_axi_rmem6___Stream2Mmap_6___mmap_RRESP;
  wire m_axi_rmem6___Stream2Mmap_6___mmap_RVALID;
  wire [511:0] m_axi_rmem6___Stream2Mmap_6___mmap_WDATA;
  wire m_axi_rmem6___Stream2Mmap_6___mmap_WLAST;
  wire m_axi_rmem6___Stream2Mmap_6___mmap_WREADY;
  wire [63:0] m_axi_rmem6___Stream2Mmap_6___mmap_WSTRB;
  wire m_axi_rmem6___Stream2Mmap_6___mmap_WVALID;
  wire [63:0] m_axi_rmem7___Mmap2Stream_7___mmap_ARADDR;
  wire [1:0] m_axi_rmem7___Mmap2Stream_7___mmap_ARBURST;
  wire [3:0] m_axi_rmem7___Mmap2Stream_7___mmap_ARCACHE;
  wire [0:0] m_axi_rmem7___Mmap2Stream_7___mmap_ARID;
  wire [7:0] m_axi_rmem7___Mmap2Stream_7___mmap_ARLEN;
  wire m_axi_rmem7___Mmap2Stream_7___mmap_ARLOCK;
  wire [2:0] m_axi_rmem7___Mmap2Stream_7___mmap_ARPROT;
  wire [3:0] m_axi_rmem7___Mmap2Stream_7___mmap_ARQOS;
  wire m_axi_rmem7___Mmap2Stream_7___mmap_ARREADY;
  wire [2:0] m_axi_rmem7___Mmap2Stream_7___mmap_ARSIZE;
  wire m_axi_rmem7___Mmap2Stream_7___mmap_ARVALID;
  wire [63:0] m_axi_rmem7___Mmap2Stream_7___mmap_AWADDR;
  wire [1:0] m_axi_rmem7___Mmap2Stream_7___mmap_AWBURST;
  wire [3:0] m_axi_rmem7___Mmap2Stream_7___mmap_AWCACHE;
  wire [0:0] m_axi_rmem7___Mmap2Stream_7___mmap_AWID;
  wire [7:0] m_axi_rmem7___Mmap2Stream_7___mmap_AWLEN;
  wire m_axi_rmem7___Mmap2Stream_7___mmap_AWLOCK;
  wire [2:0] m_axi_rmem7___Mmap2Stream_7___mmap_AWPROT;
  wire [3:0] m_axi_rmem7___Mmap2Stream_7___mmap_AWQOS;
  wire m_axi_rmem7___Mmap2Stream_7___mmap_AWREADY;
  wire [2:0] m_axi_rmem7___Mmap2Stream_7___mmap_AWSIZE;
  wire m_axi_rmem7___Mmap2Stream_7___mmap_AWVALID;
  wire [0:0] m_axi_rmem7___Mmap2Stream_7___mmap_BID;
  wire m_axi_rmem7___Mmap2Stream_7___mmap_BREADY;
  wire [1:0] m_axi_rmem7___Mmap2Stream_7___mmap_BRESP;
  wire m_axi_rmem7___Mmap2Stream_7___mmap_BVALID;
  wire [511:0] m_axi_rmem7___Mmap2Stream_7___mmap_RDATA;
  wire [0:0] m_axi_rmem7___Mmap2Stream_7___mmap_RID;
  wire m_axi_rmem7___Mmap2Stream_7___mmap_RLAST;
  wire m_axi_rmem7___Mmap2Stream_7___mmap_RREADY;
  wire [1:0] m_axi_rmem7___Mmap2Stream_7___mmap_RRESP;
  wire m_axi_rmem7___Mmap2Stream_7___mmap_RVALID;
  wire [511:0] m_axi_rmem7___Mmap2Stream_7___mmap_WDATA;
  wire m_axi_rmem7___Mmap2Stream_7___mmap_WLAST;
  wire m_axi_rmem7___Mmap2Stream_7___mmap_WREADY;
  wire [63:0] m_axi_rmem7___Mmap2Stream_7___mmap_WSTRB;
  wire m_axi_rmem7___Mmap2Stream_7___mmap_WVALID;
  wire [63:0] m_axi_rmem7___Stream2Mmap_7___mmap_ARADDR;
  wire [1:0] m_axi_rmem7___Stream2Mmap_7___mmap_ARBURST;
  wire [3:0] m_axi_rmem7___Stream2Mmap_7___mmap_ARCACHE;
  wire [0:0] m_axi_rmem7___Stream2Mmap_7___mmap_ARID;
  wire [7:0] m_axi_rmem7___Stream2Mmap_7___mmap_ARLEN;
  wire m_axi_rmem7___Stream2Mmap_7___mmap_ARLOCK;
  wire [2:0] m_axi_rmem7___Stream2Mmap_7___mmap_ARPROT;
  wire [3:0] m_axi_rmem7___Stream2Mmap_7___mmap_ARQOS;
  wire m_axi_rmem7___Stream2Mmap_7___mmap_ARREADY;
  wire [2:0] m_axi_rmem7___Stream2Mmap_7___mmap_ARSIZE;
  wire m_axi_rmem7___Stream2Mmap_7___mmap_ARVALID;
  wire [63:0] m_axi_rmem7___Stream2Mmap_7___mmap_AWADDR;
  wire [1:0] m_axi_rmem7___Stream2Mmap_7___mmap_AWBURST;
  wire [3:0] m_axi_rmem7___Stream2Mmap_7___mmap_AWCACHE;
  wire [0:0] m_axi_rmem7___Stream2Mmap_7___mmap_AWID;
  wire [7:0] m_axi_rmem7___Stream2Mmap_7___mmap_AWLEN;
  wire m_axi_rmem7___Stream2Mmap_7___mmap_AWLOCK;
  wire [2:0] m_axi_rmem7___Stream2Mmap_7___mmap_AWPROT;
  wire [3:0] m_axi_rmem7___Stream2Mmap_7___mmap_AWQOS;
  wire m_axi_rmem7___Stream2Mmap_7___mmap_AWREADY;
  wire [2:0] m_axi_rmem7___Stream2Mmap_7___mmap_AWSIZE;
  wire m_axi_rmem7___Stream2Mmap_7___mmap_AWVALID;
  wire [0:0] m_axi_rmem7___Stream2Mmap_7___mmap_BID;
  wire m_axi_rmem7___Stream2Mmap_7___mmap_BREADY;
  wire [1:0] m_axi_rmem7___Stream2Mmap_7___mmap_BRESP;
  wire m_axi_rmem7___Stream2Mmap_7___mmap_BVALID;
  wire [511:0] m_axi_rmem7___Stream2Mmap_7___mmap_RDATA;
  wire [0:0] m_axi_rmem7___Stream2Mmap_7___mmap_RID;
  wire m_axi_rmem7___Stream2Mmap_7___mmap_RLAST;
  wire m_axi_rmem7___Stream2Mmap_7___mmap_RREADY;
  wire [1:0] m_axi_rmem7___Stream2Mmap_7___mmap_RRESP;
  wire m_axi_rmem7___Stream2Mmap_7___mmap_RVALID;
  wire [511:0] m_axi_rmem7___Stream2Mmap_7___mmap_WDATA;
  wire m_axi_rmem7___Stream2Mmap_7___mmap_WLAST;
  wire m_axi_rmem7___Stream2Mmap_7___mmap_WREADY;
  wire [63:0] m_axi_rmem7___Stream2Mmap_7___mmap_WSTRB;
  wire m_axi_rmem7___Stream2Mmap_7___mmap_WVALID;
  wire [63:0] m_axi_rmem8___Mmap2Stream_8___mmap_ARADDR;
  wire [1:0] m_axi_rmem8___Mmap2Stream_8___mmap_ARBURST;
  wire [3:0] m_axi_rmem8___Mmap2Stream_8___mmap_ARCACHE;
  wire [0:0] m_axi_rmem8___Mmap2Stream_8___mmap_ARID;
  wire [7:0] m_axi_rmem8___Mmap2Stream_8___mmap_ARLEN;
  wire m_axi_rmem8___Mmap2Stream_8___mmap_ARLOCK;
  wire [2:0] m_axi_rmem8___Mmap2Stream_8___mmap_ARPROT;
  wire [3:0] m_axi_rmem8___Mmap2Stream_8___mmap_ARQOS;
  wire m_axi_rmem8___Mmap2Stream_8___mmap_ARREADY;
  wire [2:0] m_axi_rmem8___Mmap2Stream_8___mmap_ARSIZE;
  wire m_axi_rmem8___Mmap2Stream_8___mmap_ARVALID;
  wire [63:0] m_axi_rmem8___Mmap2Stream_8___mmap_AWADDR;
  wire [1:0] m_axi_rmem8___Mmap2Stream_8___mmap_AWBURST;
  wire [3:0] m_axi_rmem8___Mmap2Stream_8___mmap_AWCACHE;
  wire [0:0] m_axi_rmem8___Mmap2Stream_8___mmap_AWID;
  wire [7:0] m_axi_rmem8___Mmap2Stream_8___mmap_AWLEN;
  wire m_axi_rmem8___Mmap2Stream_8___mmap_AWLOCK;
  wire [2:0] m_axi_rmem8___Mmap2Stream_8___mmap_AWPROT;
  wire [3:0] m_axi_rmem8___Mmap2Stream_8___mmap_AWQOS;
  wire m_axi_rmem8___Mmap2Stream_8___mmap_AWREADY;
  wire [2:0] m_axi_rmem8___Mmap2Stream_8___mmap_AWSIZE;
  wire m_axi_rmem8___Mmap2Stream_8___mmap_AWVALID;
  wire [0:0] m_axi_rmem8___Mmap2Stream_8___mmap_BID;
  wire m_axi_rmem8___Mmap2Stream_8___mmap_BREADY;
  wire [1:0] m_axi_rmem8___Mmap2Stream_8___mmap_BRESP;
  wire m_axi_rmem8___Mmap2Stream_8___mmap_BVALID;
  wire [511:0] m_axi_rmem8___Mmap2Stream_8___mmap_RDATA;
  wire [0:0] m_axi_rmem8___Mmap2Stream_8___mmap_RID;
  wire m_axi_rmem8___Mmap2Stream_8___mmap_RLAST;
  wire m_axi_rmem8___Mmap2Stream_8___mmap_RREADY;
  wire [1:0] m_axi_rmem8___Mmap2Stream_8___mmap_RRESP;
  wire m_axi_rmem8___Mmap2Stream_8___mmap_RVALID;
  wire [511:0] m_axi_rmem8___Mmap2Stream_8___mmap_WDATA;
  wire m_axi_rmem8___Mmap2Stream_8___mmap_WLAST;
  wire m_axi_rmem8___Mmap2Stream_8___mmap_WREADY;
  wire [63:0] m_axi_rmem8___Mmap2Stream_8___mmap_WSTRB;
  wire m_axi_rmem8___Mmap2Stream_8___mmap_WVALID;
  wire [63:0] m_axi_rmem8___Stream2Mmap_8___mmap_ARADDR;
  wire [1:0] m_axi_rmem8___Stream2Mmap_8___mmap_ARBURST;
  wire [3:0] m_axi_rmem8___Stream2Mmap_8___mmap_ARCACHE;
  wire [0:0] m_axi_rmem8___Stream2Mmap_8___mmap_ARID;
  wire [7:0] m_axi_rmem8___Stream2Mmap_8___mmap_ARLEN;
  wire m_axi_rmem8___Stream2Mmap_8___mmap_ARLOCK;
  wire [2:0] m_axi_rmem8___Stream2Mmap_8___mmap_ARPROT;
  wire [3:0] m_axi_rmem8___Stream2Mmap_8___mmap_ARQOS;
  wire m_axi_rmem8___Stream2Mmap_8___mmap_ARREADY;
  wire [2:0] m_axi_rmem8___Stream2Mmap_8___mmap_ARSIZE;
  wire m_axi_rmem8___Stream2Mmap_8___mmap_ARVALID;
  wire [63:0] m_axi_rmem8___Stream2Mmap_8___mmap_AWADDR;
  wire [1:0] m_axi_rmem8___Stream2Mmap_8___mmap_AWBURST;
  wire [3:0] m_axi_rmem8___Stream2Mmap_8___mmap_AWCACHE;
  wire [0:0] m_axi_rmem8___Stream2Mmap_8___mmap_AWID;
  wire [7:0] m_axi_rmem8___Stream2Mmap_8___mmap_AWLEN;
  wire m_axi_rmem8___Stream2Mmap_8___mmap_AWLOCK;
  wire [2:0] m_axi_rmem8___Stream2Mmap_8___mmap_AWPROT;
  wire [3:0] m_axi_rmem8___Stream2Mmap_8___mmap_AWQOS;
  wire m_axi_rmem8___Stream2Mmap_8___mmap_AWREADY;
  wire [2:0] m_axi_rmem8___Stream2Mmap_8___mmap_AWSIZE;
  wire m_axi_rmem8___Stream2Mmap_8___mmap_AWVALID;
  wire [0:0] m_axi_rmem8___Stream2Mmap_8___mmap_BID;
  wire m_axi_rmem8___Stream2Mmap_8___mmap_BREADY;
  wire [1:0] m_axi_rmem8___Stream2Mmap_8___mmap_BRESP;
  wire m_axi_rmem8___Stream2Mmap_8___mmap_BVALID;
  wire [511:0] m_axi_rmem8___Stream2Mmap_8___mmap_RDATA;
  wire [0:0] m_axi_rmem8___Stream2Mmap_8___mmap_RID;
  wire m_axi_rmem8___Stream2Mmap_8___mmap_RLAST;
  wire m_axi_rmem8___Stream2Mmap_8___mmap_RREADY;
  wire [1:0] m_axi_rmem8___Stream2Mmap_8___mmap_RRESP;
  wire m_axi_rmem8___Stream2Mmap_8___mmap_RVALID;
  wire [511:0] m_axi_rmem8___Stream2Mmap_8___mmap_WDATA;
  wire m_axi_rmem8___Stream2Mmap_8___mmap_WLAST;
  wire m_axi_rmem8___Stream2Mmap_8___mmap_WREADY;
  wire [63:0] m_axi_rmem8___Stream2Mmap_8___mmap_WSTRB;
  wire m_axi_rmem8___Stream2Mmap_8___mmap_WVALID;
  wire [63:0] m_axi_rmem9___Mmap2Stream_9___mmap_ARADDR;
  wire [1:0] m_axi_rmem9___Mmap2Stream_9___mmap_ARBURST;
  wire [3:0] m_axi_rmem9___Mmap2Stream_9___mmap_ARCACHE;
  wire [0:0] m_axi_rmem9___Mmap2Stream_9___mmap_ARID;
  wire [7:0] m_axi_rmem9___Mmap2Stream_9___mmap_ARLEN;
  wire m_axi_rmem9___Mmap2Stream_9___mmap_ARLOCK;
  wire [2:0] m_axi_rmem9___Mmap2Stream_9___mmap_ARPROT;
  wire [3:0] m_axi_rmem9___Mmap2Stream_9___mmap_ARQOS;
  wire m_axi_rmem9___Mmap2Stream_9___mmap_ARREADY;
  wire [2:0] m_axi_rmem9___Mmap2Stream_9___mmap_ARSIZE;
  wire m_axi_rmem9___Mmap2Stream_9___mmap_ARVALID;
  wire [63:0] m_axi_rmem9___Mmap2Stream_9___mmap_AWADDR;
  wire [1:0] m_axi_rmem9___Mmap2Stream_9___mmap_AWBURST;
  wire [3:0] m_axi_rmem9___Mmap2Stream_9___mmap_AWCACHE;
  wire [0:0] m_axi_rmem9___Mmap2Stream_9___mmap_AWID;
  wire [7:0] m_axi_rmem9___Mmap2Stream_9___mmap_AWLEN;
  wire m_axi_rmem9___Mmap2Stream_9___mmap_AWLOCK;
  wire [2:0] m_axi_rmem9___Mmap2Stream_9___mmap_AWPROT;
  wire [3:0] m_axi_rmem9___Mmap2Stream_9___mmap_AWQOS;
  wire m_axi_rmem9___Mmap2Stream_9___mmap_AWREADY;
  wire [2:0] m_axi_rmem9___Mmap2Stream_9___mmap_AWSIZE;
  wire m_axi_rmem9___Mmap2Stream_9___mmap_AWVALID;
  wire [0:0] m_axi_rmem9___Mmap2Stream_9___mmap_BID;
  wire m_axi_rmem9___Mmap2Stream_9___mmap_BREADY;
  wire [1:0] m_axi_rmem9___Mmap2Stream_9___mmap_BRESP;
  wire m_axi_rmem9___Mmap2Stream_9___mmap_BVALID;
  wire [511:0] m_axi_rmem9___Mmap2Stream_9___mmap_RDATA;
  wire [0:0] m_axi_rmem9___Mmap2Stream_9___mmap_RID;
  wire m_axi_rmem9___Mmap2Stream_9___mmap_RLAST;
  wire m_axi_rmem9___Mmap2Stream_9___mmap_RREADY;
  wire [1:0] m_axi_rmem9___Mmap2Stream_9___mmap_RRESP;
  wire m_axi_rmem9___Mmap2Stream_9___mmap_RVALID;
  wire [511:0] m_axi_rmem9___Mmap2Stream_9___mmap_WDATA;
  wire m_axi_rmem9___Mmap2Stream_9___mmap_WLAST;
  wire m_axi_rmem9___Mmap2Stream_9___mmap_WREADY;
  wire [63:0] m_axi_rmem9___Mmap2Stream_9___mmap_WSTRB;
  wire m_axi_rmem9___Mmap2Stream_9___mmap_WVALID;
  wire [63:0] m_axi_rmem9___Stream2Mmap_9___mmap_ARADDR;
  wire [1:0] m_axi_rmem9___Stream2Mmap_9___mmap_ARBURST;
  wire [3:0] m_axi_rmem9___Stream2Mmap_9___mmap_ARCACHE;
  wire [0:0] m_axi_rmem9___Stream2Mmap_9___mmap_ARID;
  wire [7:0] m_axi_rmem9___Stream2Mmap_9___mmap_ARLEN;
  wire m_axi_rmem9___Stream2Mmap_9___mmap_ARLOCK;
  wire [2:0] m_axi_rmem9___Stream2Mmap_9___mmap_ARPROT;
  wire [3:0] m_axi_rmem9___Stream2Mmap_9___mmap_ARQOS;
  wire m_axi_rmem9___Stream2Mmap_9___mmap_ARREADY;
  wire [2:0] m_axi_rmem9___Stream2Mmap_9___mmap_ARSIZE;
  wire m_axi_rmem9___Stream2Mmap_9___mmap_ARVALID;
  wire [63:0] m_axi_rmem9___Stream2Mmap_9___mmap_AWADDR;
  wire [1:0] m_axi_rmem9___Stream2Mmap_9___mmap_AWBURST;
  wire [3:0] m_axi_rmem9___Stream2Mmap_9___mmap_AWCACHE;
  wire [0:0] m_axi_rmem9___Stream2Mmap_9___mmap_AWID;
  wire [7:0] m_axi_rmem9___Stream2Mmap_9___mmap_AWLEN;
  wire m_axi_rmem9___Stream2Mmap_9___mmap_AWLOCK;
  wire [2:0] m_axi_rmem9___Stream2Mmap_9___mmap_AWPROT;
  wire [3:0] m_axi_rmem9___Stream2Mmap_9___mmap_AWQOS;
  wire m_axi_rmem9___Stream2Mmap_9___mmap_AWREADY;
  wire [2:0] m_axi_rmem9___Stream2Mmap_9___mmap_AWSIZE;
  wire m_axi_rmem9___Stream2Mmap_9___mmap_AWVALID;
  wire [0:0] m_axi_rmem9___Stream2Mmap_9___mmap_BID;
  wire m_axi_rmem9___Stream2Mmap_9___mmap_BREADY;
  wire [1:0] m_axi_rmem9___Stream2Mmap_9___mmap_BRESP;
  wire m_axi_rmem9___Stream2Mmap_9___mmap_BVALID;
  wire [511:0] m_axi_rmem9___Stream2Mmap_9___mmap_RDATA;
  wire [0:0] m_axi_rmem9___Stream2Mmap_9___mmap_RID;
  wire m_axi_rmem9___Stream2Mmap_9___mmap_RLAST;
  wire m_axi_rmem9___Stream2Mmap_9___mmap_RREADY;
  wire [1:0] m_axi_rmem9___Stream2Mmap_9___mmap_RRESP;
  wire m_axi_rmem9___Stream2Mmap_9___mmap_RVALID;
  wire [511:0] m_axi_rmem9___Stream2Mmap_9___mmap_WDATA;
  wire m_axi_rmem9___Stream2Mmap_9___mmap_WLAST;
  wire m_axi_rmem9___Stream2Mmap_9___mmap_WREADY;
  wire [63:0] m_axi_rmem9___Stream2Mmap_9___mmap_WSTRB;
  wire m_axi_rmem9___Stream2Mmap_9___mmap_WVALID;
  wire [63:0] m_axi_rmem10___Mmap2Stream_10___mmap_ARADDR;
  wire [1:0] m_axi_rmem10___Mmap2Stream_10___mmap_ARBURST;
  wire [3:0] m_axi_rmem10___Mmap2Stream_10___mmap_ARCACHE;
  wire [0:0] m_axi_rmem10___Mmap2Stream_10___mmap_ARID;
  wire [7:0] m_axi_rmem10___Mmap2Stream_10___mmap_ARLEN;
  wire m_axi_rmem10___Mmap2Stream_10___mmap_ARLOCK;
  wire [2:0] m_axi_rmem10___Mmap2Stream_10___mmap_ARPROT;
  wire [3:0] m_axi_rmem10___Mmap2Stream_10___mmap_ARQOS;
  wire m_axi_rmem10___Mmap2Stream_10___mmap_ARREADY;
  wire [2:0] m_axi_rmem10___Mmap2Stream_10___mmap_ARSIZE;
  wire m_axi_rmem10___Mmap2Stream_10___mmap_ARVALID;
  wire [63:0] m_axi_rmem10___Mmap2Stream_10___mmap_AWADDR;
  wire [1:0] m_axi_rmem10___Mmap2Stream_10___mmap_AWBURST;
  wire [3:0] m_axi_rmem10___Mmap2Stream_10___mmap_AWCACHE;
  wire [0:0] m_axi_rmem10___Mmap2Stream_10___mmap_AWID;
  wire [7:0] m_axi_rmem10___Mmap2Stream_10___mmap_AWLEN;
  wire m_axi_rmem10___Mmap2Stream_10___mmap_AWLOCK;
  wire [2:0] m_axi_rmem10___Mmap2Stream_10___mmap_AWPROT;
  wire [3:0] m_axi_rmem10___Mmap2Stream_10___mmap_AWQOS;
  wire m_axi_rmem10___Mmap2Stream_10___mmap_AWREADY;
  wire [2:0] m_axi_rmem10___Mmap2Stream_10___mmap_AWSIZE;
  wire m_axi_rmem10___Mmap2Stream_10___mmap_AWVALID;
  wire [0:0] m_axi_rmem10___Mmap2Stream_10___mmap_BID;
  wire m_axi_rmem10___Mmap2Stream_10___mmap_BREADY;
  wire [1:0] m_axi_rmem10___Mmap2Stream_10___mmap_BRESP;
  wire m_axi_rmem10___Mmap2Stream_10___mmap_BVALID;
  wire [511:0] m_axi_rmem10___Mmap2Stream_10___mmap_RDATA;
  wire [0:0] m_axi_rmem10___Mmap2Stream_10___mmap_RID;
  wire m_axi_rmem10___Mmap2Stream_10___mmap_RLAST;
  wire m_axi_rmem10___Mmap2Stream_10___mmap_RREADY;
  wire [1:0] m_axi_rmem10___Mmap2Stream_10___mmap_RRESP;
  wire m_axi_rmem10___Mmap2Stream_10___mmap_RVALID;
  wire [511:0] m_axi_rmem10___Mmap2Stream_10___mmap_WDATA;
  wire m_axi_rmem10___Mmap2Stream_10___mmap_WLAST;
  wire m_axi_rmem10___Mmap2Stream_10___mmap_WREADY;
  wire [63:0] m_axi_rmem10___Mmap2Stream_10___mmap_WSTRB;
  wire m_axi_rmem10___Mmap2Stream_10___mmap_WVALID;
  wire [63:0] m_axi_rmem10___Stream2Mmap_10___mmap_ARADDR;
  wire [1:0] m_axi_rmem10___Stream2Mmap_10___mmap_ARBURST;
  wire [3:0] m_axi_rmem10___Stream2Mmap_10___mmap_ARCACHE;
  wire [0:0] m_axi_rmem10___Stream2Mmap_10___mmap_ARID;
  wire [7:0] m_axi_rmem10___Stream2Mmap_10___mmap_ARLEN;
  wire m_axi_rmem10___Stream2Mmap_10___mmap_ARLOCK;
  wire [2:0] m_axi_rmem10___Stream2Mmap_10___mmap_ARPROT;
  wire [3:0] m_axi_rmem10___Stream2Mmap_10___mmap_ARQOS;
  wire m_axi_rmem10___Stream2Mmap_10___mmap_ARREADY;
  wire [2:0] m_axi_rmem10___Stream2Mmap_10___mmap_ARSIZE;
  wire m_axi_rmem10___Stream2Mmap_10___mmap_ARVALID;
  wire [63:0] m_axi_rmem10___Stream2Mmap_10___mmap_AWADDR;
  wire [1:0] m_axi_rmem10___Stream2Mmap_10___mmap_AWBURST;
  wire [3:0] m_axi_rmem10___Stream2Mmap_10___mmap_AWCACHE;
  wire [0:0] m_axi_rmem10___Stream2Mmap_10___mmap_AWID;
  wire [7:0] m_axi_rmem10___Stream2Mmap_10___mmap_AWLEN;
  wire m_axi_rmem10___Stream2Mmap_10___mmap_AWLOCK;
  wire [2:0] m_axi_rmem10___Stream2Mmap_10___mmap_AWPROT;
  wire [3:0] m_axi_rmem10___Stream2Mmap_10___mmap_AWQOS;
  wire m_axi_rmem10___Stream2Mmap_10___mmap_AWREADY;
  wire [2:0] m_axi_rmem10___Stream2Mmap_10___mmap_AWSIZE;
  wire m_axi_rmem10___Stream2Mmap_10___mmap_AWVALID;
  wire [0:0] m_axi_rmem10___Stream2Mmap_10___mmap_BID;
  wire m_axi_rmem10___Stream2Mmap_10___mmap_BREADY;
  wire [1:0] m_axi_rmem10___Stream2Mmap_10___mmap_BRESP;
  wire m_axi_rmem10___Stream2Mmap_10___mmap_BVALID;
  wire [511:0] m_axi_rmem10___Stream2Mmap_10___mmap_RDATA;
  wire [0:0] m_axi_rmem10___Stream2Mmap_10___mmap_RID;
  wire m_axi_rmem10___Stream2Mmap_10___mmap_RLAST;
  wire m_axi_rmem10___Stream2Mmap_10___mmap_RREADY;
  wire [1:0] m_axi_rmem10___Stream2Mmap_10___mmap_RRESP;
  wire m_axi_rmem10___Stream2Mmap_10___mmap_RVALID;
  wire [511:0] m_axi_rmem10___Stream2Mmap_10___mmap_WDATA;
  wire m_axi_rmem10___Stream2Mmap_10___mmap_WLAST;
  wire m_axi_rmem10___Stream2Mmap_10___mmap_WREADY;
  wire [63:0] m_axi_rmem10___Stream2Mmap_10___mmap_WSTRB;
  wire m_axi_rmem10___Stream2Mmap_10___mmap_WVALID;
  wire [63:0] m_axi_rmem11___Mmap2Stream_11___mmap_ARADDR;
  wire [1:0] m_axi_rmem11___Mmap2Stream_11___mmap_ARBURST;
  wire [3:0] m_axi_rmem11___Mmap2Stream_11___mmap_ARCACHE;
  wire [0:0] m_axi_rmem11___Mmap2Stream_11___mmap_ARID;
  wire [7:0] m_axi_rmem11___Mmap2Stream_11___mmap_ARLEN;
  wire m_axi_rmem11___Mmap2Stream_11___mmap_ARLOCK;
  wire [2:0] m_axi_rmem11___Mmap2Stream_11___mmap_ARPROT;
  wire [3:0] m_axi_rmem11___Mmap2Stream_11___mmap_ARQOS;
  wire m_axi_rmem11___Mmap2Stream_11___mmap_ARREADY;
  wire [2:0] m_axi_rmem11___Mmap2Stream_11___mmap_ARSIZE;
  wire m_axi_rmem11___Mmap2Stream_11___mmap_ARVALID;
  wire [63:0] m_axi_rmem11___Mmap2Stream_11___mmap_AWADDR;
  wire [1:0] m_axi_rmem11___Mmap2Stream_11___mmap_AWBURST;
  wire [3:0] m_axi_rmem11___Mmap2Stream_11___mmap_AWCACHE;
  wire [0:0] m_axi_rmem11___Mmap2Stream_11___mmap_AWID;
  wire [7:0] m_axi_rmem11___Mmap2Stream_11___mmap_AWLEN;
  wire m_axi_rmem11___Mmap2Stream_11___mmap_AWLOCK;
  wire [2:0] m_axi_rmem11___Mmap2Stream_11___mmap_AWPROT;
  wire [3:0] m_axi_rmem11___Mmap2Stream_11___mmap_AWQOS;
  wire m_axi_rmem11___Mmap2Stream_11___mmap_AWREADY;
  wire [2:0] m_axi_rmem11___Mmap2Stream_11___mmap_AWSIZE;
  wire m_axi_rmem11___Mmap2Stream_11___mmap_AWVALID;
  wire [0:0] m_axi_rmem11___Mmap2Stream_11___mmap_BID;
  wire m_axi_rmem11___Mmap2Stream_11___mmap_BREADY;
  wire [1:0] m_axi_rmem11___Mmap2Stream_11___mmap_BRESP;
  wire m_axi_rmem11___Mmap2Stream_11___mmap_BVALID;
  wire [511:0] m_axi_rmem11___Mmap2Stream_11___mmap_RDATA;
  wire [0:0] m_axi_rmem11___Mmap2Stream_11___mmap_RID;
  wire m_axi_rmem11___Mmap2Stream_11___mmap_RLAST;
  wire m_axi_rmem11___Mmap2Stream_11___mmap_RREADY;
  wire [1:0] m_axi_rmem11___Mmap2Stream_11___mmap_RRESP;
  wire m_axi_rmem11___Mmap2Stream_11___mmap_RVALID;
  wire [511:0] m_axi_rmem11___Mmap2Stream_11___mmap_WDATA;
  wire m_axi_rmem11___Mmap2Stream_11___mmap_WLAST;
  wire m_axi_rmem11___Mmap2Stream_11___mmap_WREADY;
  wire [63:0] m_axi_rmem11___Mmap2Stream_11___mmap_WSTRB;
  wire m_axi_rmem11___Mmap2Stream_11___mmap_WVALID;
  wire [63:0] m_axi_rmem11___Stream2Mmap_11___mmap_ARADDR;
  wire [1:0] m_axi_rmem11___Stream2Mmap_11___mmap_ARBURST;
  wire [3:0] m_axi_rmem11___Stream2Mmap_11___mmap_ARCACHE;
  wire [0:0] m_axi_rmem11___Stream2Mmap_11___mmap_ARID;
  wire [7:0] m_axi_rmem11___Stream2Mmap_11___mmap_ARLEN;
  wire m_axi_rmem11___Stream2Mmap_11___mmap_ARLOCK;
  wire [2:0] m_axi_rmem11___Stream2Mmap_11___mmap_ARPROT;
  wire [3:0] m_axi_rmem11___Stream2Mmap_11___mmap_ARQOS;
  wire m_axi_rmem11___Stream2Mmap_11___mmap_ARREADY;
  wire [2:0] m_axi_rmem11___Stream2Mmap_11___mmap_ARSIZE;
  wire m_axi_rmem11___Stream2Mmap_11___mmap_ARVALID;
  wire [63:0] m_axi_rmem11___Stream2Mmap_11___mmap_AWADDR;
  wire [1:0] m_axi_rmem11___Stream2Mmap_11___mmap_AWBURST;
  wire [3:0] m_axi_rmem11___Stream2Mmap_11___mmap_AWCACHE;
  wire [0:0] m_axi_rmem11___Stream2Mmap_11___mmap_AWID;
  wire [7:0] m_axi_rmem11___Stream2Mmap_11___mmap_AWLEN;
  wire m_axi_rmem11___Stream2Mmap_11___mmap_AWLOCK;
  wire [2:0] m_axi_rmem11___Stream2Mmap_11___mmap_AWPROT;
  wire [3:0] m_axi_rmem11___Stream2Mmap_11___mmap_AWQOS;
  wire m_axi_rmem11___Stream2Mmap_11___mmap_AWREADY;
  wire [2:0] m_axi_rmem11___Stream2Mmap_11___mmap_AWSIZE;
  wire m_axi_rmem11___Stream2Mmap_11___mmap_AWVALID;
  wire [0:0] m_axi_rmem11___Stream2Mmap_11___mmap_BID;
  wire m_axi_rmem11___Stream2Mmap_11___mmap_BREADY;
  wire [1:0] m_axi_rmem11___Stream2Mmap_11___mmap_BRESP;
  wire m_axi_rmem11___Stream2Mmap_11___mmap_BVALID;
  wire [511:0] m_axi_rmem11___Stream2Mmap_11___mmap_RDATA;
  wire [0:0] m_axi_rmem11___Stream2Mmap_11___mmap_RID;
  wire m_axi_rmem11___Stream2Mmap_11___mmap_RLAST;
  wire m_axi_rmem11___Stream2Mmap_11___mmap_RREADY;
  wire [1:0] m_axi_rmem11___Stream2Mmap_11___mmap_RRESP;
  wire m_axi_rmem11___Stream2Mmap_11___mmap_RVALID;
  wire [511:0] m_axi_rmem11___Stream2Mmap_11___mmap_WDATA;
  wire m_axi_rmem11___Stream2Mmap_11___mmap_WLAST;
  wire m_axi_rmem11___Stream2Mmap_11___mmap_WREADY;
  wire [63:0] m_axi_rmem11___Stream2Mmap_11___mmap_WSTRB;
  wire m_axi_rmem11___Stream2Mmap_11___mmap_WVALID;
  wire [63:0] m_axi_rmem12___Mmap2Stream_12___mmap_ARADDR;
  wire [1:0] m_axi_rmem12___Mmap2Stream_12___mmap_ARBURST;
  wire [3:0] m_axi_rmem12___Mmap2Stream_12___mmap_ARCACHE;
  wire [0:0] m_axi_rmem12___Mmap2Stream_12___mmap_ARID;
  wire [7:0] m_axi_rmem12___Mmap2Stream_12___mmap_ARLEN;
  wire m_axi_rmem12___Mmap2Stream_12___mmap_ARLOCK;
  wire [2:0] m_axi_rmem12___Mmap2Stream_12___mmap_ARPROT;
  wire [3:0] m_axi_rmem12___Mmap2Stream_12___mmap_ARQOS;
  wire m_axi_rmem12___Mmap2Stream_12___mmap_ARREADY;
  wire [2:0] m_axi_rmem12___Mmap2Stream_12___mmap_ARSIZE;
  wire m_axi_rmem12___Mmap2Stream_12___mmap_ARVALID;
  wire [63:0] m_axi_rmem12___Mmap2Stream_12___mmap_AWADDR;
  wire [1:0] m_axi_rmem12___Mmap2Stream_12___mmap_AWBURST;
  wire [3:0] m_axi_rmem12___Mmap2Stream_12___mmap_AWCACHE;
  wire [0:0] m_axi_rmem12___Mmap2Stream_12___mmap_AWID;
  wire [7:0] m_axi_rmem12___Mmap2Stream_12___mmap_AWLEN;
  wire m_axi_rmem12___Mmap2Stream_12___mmap_AWLOCK;
  wire [2:0] m_axi_rmem12___Mmap2Stream_12___mmap_AWPROT;
  wire [3:0] m_axi_rmem12___Mmap2Stream_12___mmap_AWQOS;
  wire m_axi_rmem12___Mmap2Stream_12___mmap_AWREADY;
  wire [2:0] m_axi_rmem12___Mmap2Stream_12___mmap_AWSIZE;
  wire m_axi_rmem12___Mmap2Stream_12___mmap_AWVALID;
  wire [0:0] m_axi_rmem12___Mmap2Stream_12___mmap_BID;
  wire m_axi_rmem12___Mmap2Stream_12___mmap_BREADY;
  wire [1:0] m_axi_rmem12___Mmap2Stream_12___mmap_BRESP;
  wire m_axi_rmem12___Mmap2Stream_12___mmap_BVALID;
  wire [511:0] m_axi_rmem12___Mmap2Stream_12___mmap_RDATA;
  wire [0:0] m_axi_rmem12___Mmap2Stream_12___mmap_RID;
  wire m_axi_rmem12___Mmap2Stream_12___mmap_RLAST;
  wire m_axi_rmem12___Mmap2Stream_12___mmap_RREADY;
  wire [1:0] m_axi_rmem12___Mmap2Stream_12___mmap_RRESP;
  wire m_axi_rmem12___Mmap2Stream_12___mmap_RVALID;
  wire [511:0] m_axi_rmem12___Mmap2Stream_12___mmap_WDATA;
  wire m_axi_rmem12___Mmap2Stream_12___mmap_WLAST;
  wire m_axi_rmem12___Mmap2Stream_12___mmap_WREADY;
  wire [63:0] m_axi_rmem12___Mmap2Stream_12___mmap_WSTRB;
  wire m_axi_rmem12___Mmap2Stream_12___mmap_WVALID;
  wire [63:0] m_axi_rmem12___Stream2Mmap_12___mmap_ARADDR;
  wire [1:0] m_axi_rmem12___Stream2Mmap_12___mmap_ARBURST;
  wire [3:0] m_axi_rmem12___Stream2Mmap_12___mmap_ARCACHE;
  wire [0:0] m_axi_rmem12___Stream2Mmap_12___mmap_ARID;
  wire [7:0] m_axi_rmem12___Stream2Mmap_12___mmap_ARLEN;
  wire m_axi_rmem12___Stream2Mmap_12___mmap_ARLOCK;
  wire [2:0] m_axi_rmem12___Stream2Mmap_12___mmap_ARPROT;
  wire [3:0] m_axi_rmem12___Stream2Mmap_12___mmap_ARQOS;
  wire m_axi_rmem12___Stream2Mmap_12___mmap_ARREADY;
  wire [2:0] m_axi_rmem12___Stream2Mmap_12___mmap_ARSIZE;
  wire m_axi_rmem12___Stream2Mmap_12___mmap_ARVALID;
  wire [63:0] m_axi_rmem12___Stream2Mmap_12___mmap_AWADDR;
  wire [1:0] m_axi_rmem12___Stream2Mmap_12___mmap_AWBURST;
  wire [3:0] m_axi_rmem12___Stream2Mmap_12___mmap_AWCACHE;
  wire [0:0] m_axi_rmem12___Stream2Mmap_12___mmap_AWID;
  wire [7:0] m_axi_rmem12___Stream2Mmap_12___mmap_AWLEN;
  wire m_axi_rmem12___Stream2Mmap_12___mmap_AWLOCK;
  wire [2:0] m_axi_rmem12___Stream2Mmap_12___mmap_AWPROT;
  wire [3:0] m_axi_rmem12___Stream2Mmap_12___mmap_AWQOS;
  wire m_axi_rmem12___Stream2Mmap_12___mmap_AWREADY;
  wire [2:0] m_axi_rmem12___Stream2Mmap_12___mmap_AWSIZE;
  wire m_axi_rmem12___Stream2Mmap_12___mmap_AWVALID;
  wire [0:0] m_axi_rmem12___Stream2Mmap_12___mmap_BID;
  wire m_axi_rmem12___Stream2Mmap_12___mmap_BREADY;
  wire [1:0] m_axi_rmem12___Stream2Mmap_12___mmap_BRESP;
  wire m_axi_rmem12___Stream2Mmap_12___mmap_BVALID;
  wire [511:0] m_axi_rmem12___Stream2Mmap_12___mmap_RDATA;
  wire [0:0] m_axi_rmem12___Stream2Mmap_12___mmap_RID;
  wire m_axi_rmem12___Stream2Mmap_12___mmap_RLAST;
  wire m_axi_rmem12___Stream2Mmap_12___mmap_RREADY;
  wire [1:0] m_axi_rmem12___Stream2Mmap_12___mmap_RRESP;
  wire m_axi_rmem12___Stream2Mmap_12___mmap_RVALID;
  wire [511:0] m_axi_rmem12___Stream2Mmap_12___mmap_WDATA;
  wire m_axi_rmem12___Stream2Mmap_12___mmap_WLAST;
  wire m_axi_rmem12___Stream2Mmap_12___mmap_WREADY;
  wire [63:0] m_axi_rmem12___Stream2Mmap_12___mmap_WSTRB;
  wire m_axi_rmem12___Stream2Mmap_12___mmap_WVALID;
  wire [63:0] m_axi_rmem13___Mmap2Stream_13___mmap_ARADDR;
  wire [1:0] m_axi_rmem13___Mmap2Stream_13___mmap_ARBURST;
  wire [3:0] m_axi_rmem13___Mmap2Stream_13___mmap_ARCACHE;
  wire [0:0] m_axi_rmem13___Mmap2Stream_13___mmap_ARID;
  wire [7:0] m_axi_rmem13___Mmap2Stream_13___mmap_ARLEN;
  wire m_axi_rmem13___Mmap2Stream_13___mmap_ARLOCK;
  wire [2:0] m_axi_rmem13___Mmap2Stream_13___mmap_ARPROT;
  wire [3:0] m_axi_rmem13___Mmap2Stream_13___mmap_ARQOS;
  wire m_axi_rmem13___Mmap2Stream_13___mmap_ARREADY;
  wire [2:0] m_axi_rmem13___Mmap2Stream_13___mmap_ARSIZE;
  wire m_axi_rmem13___Mmap2Stream_13___mmap_ARVALID;
  wire [63:0] m_axi_rmem13___Mmap2Stream_13___mmap_AWADDR;
  wire [1:0] m_axi_rmem13___Mmap2Stream_13___mmap_AWBURST;
  wire [3:0] m_axi_rmem13___Mmap2Stream_13___mmap_AWCACHE;
  wire [0:0] m_axi_rmem13___Mmap2Stream_13___mmap_AWID;
  wire [7:0] m_axi_rmem13___Mmap2Stream_13___mmap_AWLEN;
  wire m_axi_rmem13___Mmap2Stream_13___mmap_AWLOCK;
  wire [2:0] m_axi_rmem13___Mmap2Stream_13___mmap_AWPROT;
  wire [3:0] m_axi_rmem13___Mmap2Stream_13___mmap_AWQOS;
  wire m_axi_rmem13___Mmap2Stream_13___mmap_AWREADY;
  wire [2:0] m_axi_rmem13___Mmap2Stream_13___mmap_AWSIZE;
  wire m_axi_rmem13___Mmap2Stream_13___mmap_AWVALID;
  wire [0:0] m_axi_rmem13___Mmap2Stream_13___mmap_BID;
  wire m_axi_rmem13___Mmap2Stream_13___mmap_BREADY;
  wire [1:0] m_axi_rmem13___Mmap2Stream_13___mmap_BRESP;
  wire m_axi_rmem13___Mmap2Stream_13___mmap_BVALID;
  wire [511:0] m_axi_rmem13___Mmap2Stream_13___mmap_RDATA;
  wire [0:0] m_axi_rmem13___Mmap2Stream_13___mmap_RID;
  wire m_axi_rmem13___Mmap2Stream_13___mmap_RLAST;
  wire m_axi_rmem13___Mmap2Stream_13___mmap_RREADY;
  wire [1:0] m_axi_rmem13___Mmap2Stream_13___mmap_RRESP;
  wire m_axi_rmem13___Mmap2Stream_13___mmap_RVALID;
  wire [511:0] m_axi_rmem13___Mmap2Stream_13___mmap_WDATA;
  wire m_axi_rmem13___Mmap2Stream_13___mmap_WLAST;
  wire m_axi_rmem13___Mmap2Stream_13___mmap_WREADY;
  wire [63:0] m_axi_rmem13___Mmap2Stream_13___mmap_WSTRB;
  wire m_axi_rmem13___Mmap2Stream_13___mmap_WVALID;
  wire [63:0] m_axi_rmem13___Stream2Mmap_13___mmap_ARADDR;
  wire [1:0] m_axi_rmem13___Stream2Mmap_13___mmap_ARBURST;
  wire [3:0] m_axi_rmem13___Stream2Mmap_13___mmap_ARCACHE;
  wire [0:0] m_axi_rmem13___Stream2Mmap_13___mmap_ARID;
  wire [7:0] m_axi_rmem13___Stream2Mmap_13___mmap_ARLEN;
  wire m_axi_rmem13___Stream2Mmap_13___mmap_ARLOCK;
  wire [2:0] m_axi_rmem13___Stream2Mmap_13___mmap_ARPROT;
  wire [3:0] m_axi_rmem13___Stream2Mmap_13___mmap_ARQOS;
  wire m_axi_rmem13___Stream2Mmap_13___mmap_ARREADY;
  wire [2:0] m_axi_rmem13___Stream2Mmap_13___mmap_ARSIZE;
  wire m_axi_rmem13___Stream2Mmap_13___mmap_ARVALID;
  wire [63:0] m_axi_rmem13___Stream2Mmap_13___mmap_AWADDR;
  wire [1:0] m_axi_rmem13___Stream2Mmap_13___mmap_AWBURST;
  wire [3:0] m_axi_rmem13___Stream2Mmap_13___mmap_AWCACHE;
  wire [0:0] m_axi_rmem13___Stream2Mmap_13___mmap_AWID;
  wire [7:0] m_axi_rmem13___Stream2Mmap_13___mmap_AWLEN;
  wire m_axi_rmem13___Stream2Mmap_13___mmap_AWLOCK;
  wire [2:0] m_axi_rmem13___Stream2Mmap_13___mmap_AWPROT;
  wire [3:0] m_axi_rmem13___Stream2Mmap_13___mmap_AWQOS;
  wire m_axi_rmem13___Stream2Mmap_13___mmap_AWREADY;
  wire [2:0] m_axi_rmem13___Stream2Mmap_13___mmap_AWSIZE;
  wire m_axi_rmem13___Stream2Mmap_13___mmap_AWVALID;
  wire [0:0] m_axi_rmem13___Stream2Mmap_13___mmap_BID;
  wire m_axi_rmem13___Stream2Mmap_13___mmap_BREADY;
  wire [1:0] m_axi_rmem13___Stream2Mmap_13___mmap_BRESP;
  wire m_axi_rmem13___Stream2Mmap_13___mmap_BVALID;
  wire [511:0] m_axi_rmem13___Stream2Mmap_13___mmap_RDATA;
  wire [0:0] m_axi_rmem13___Stream2Mmap_13___mmap_RID;
  wire m_axi_rmem13___Stream2Mmap_13___mmap_RLAST;
  wire m_axi_rmem13___Stream2Mmap_13___mmap_RREADY;
  wire [1:0] m_axi_rmem13___Stream2Mmap_13___mmap_RRESP;
  wire m_axi_rmem13___Stream2Mmap_13___mmap_RVALID;
  wire [511:0] m_axi_rmem13___Stream2Mmap_13___mmap_WDATA;
  wire m_axi_rmem13___Stream2Mmap_13___mmap_WLAST;
  wire m_axi_rmem13___Stream2Mmap_13___mmap_WREADY;
  wire [63:0] m_axi_rmem13___Stream2Mmap_13___mmap_WSTRB;
  wire m_axi_rmem13___Stream2Mmap_13___mmap_WVALID;
  wire [63:0] m_axi_rmem14___Mmap2Stream_14___mmap_ARADDR;
  wire [1:0] m_axi_rmem14___Mmap2Stream_14___mmap_ARBURST;
  wire [3:0] m_axi_rmem14___Mmap2Stream_14___mmap_ARCACHE;
  wire [0:0] m_axi_rmem14___Mmap2Stream_14___mmap_ARID;
  wire [7:0] m_axi_rmem14___Mmap2Stream_14___mmap_ARLEN;
  wire m_axi_rmem14___Mmap2Stream_14___mmap_ARLOCK;
  wire [2:0] m_axi_rmem14___Mmap2Stream_14___mmap_ARPROT;
  wire [3:0] m_axi_rmem14___Mmap2Stream_14___mmap_ARQOS;
  wire m_axi_rmem14___Mmap2Stream_14___mmap_ARREADY;
  wire [2:0] m_axi_rmem14___Mmap2Stream_14___mmap_ARSIZE;
  wire m_axi_rmem14___Mmap2Stream_14___mmap_ARVALID;
  wire [63:0] m_axi_rmem14___Mmap2Stream_14___mmap_AWADDR;
  wire [1:0] m_axi_rmem14___Mmap2Stream_14___mmap_AWBURST;
  wire [3:0] m_axi_rmem14___Mmap2Stream_14___mmap_AWCACHE;
  wire [0:0] m_axi_rmem14___Mmap2Stream_14___mmap_AWID;
  wire [7:0] m_axi_rmem14___Mmap2Stream_14___mmap_AWLEN;
  wire m_axi_rmem14___Mmap2Stream_14___mmap_AWLOCK;
  wire [2:0] m_axi_rmem14___Mmap2Stream_14___mmap_AWPROT;
  wire [3:0] m_axi_rmem14___Mmap2Stream_14___mmap_AWQOS;
  wire m_axi_rmem14___Mmap2Stream_14___mmap_AWREADY;
  wire [2:0] m_axi_rmem14___Mmap2Stream_14___mmap_AWSIZE;
  wire m_axi_rmem14___Mmap2Stream_14___mmap_AWVALID;
  wire [0:0] m_axi_rmem14___Mmap2Stream_14___mmap_BID;
  wire m_axi_rmem14___Mmap2Stream_14___mmap_BREADY;
  wire [1:0] m_axi_rmem14___Mmap2Stream_14___mmap_BRESP;
  wire m_axi_rmem14___Mmap2Stream_14___mmap_BVALID;
  wire [511:0] m_axi_rmem14___Mmap2Stream_14___mmap_RDATA;
  wire [0:0] m_axi_rmem14___Mmap2Stream_14___mmap_RID;
  wire m_axi_rmem14___Mmap2Stream_14___mmap_RLAST;
  wire m_axi_rmem14___Mmap2Stream_14___mmap_RREADY;
  wire [1:0] m_axi_rmem14___Mmap2Stream_14___mmap_RRESP;
  wire m_axi_rmem14___Mmap2Stream_14___mmap_RVALID;
  wire [511:0] m_axi_rmem14___Mmap2Stream_14___mmap_WDATA;
  wire m_axi_rmem14___Mmap2Stream_14___mmap_WLAST;
  wire m_axi_rmem14___Mmap2Stream_14___mmap_WREADY;
  wire [63:0] m_axi_rmem14___Mmap2Stream_14___mmap_WSTRB;
  wire m_axi_rmem14___Mmap2Stream_14___mmap_WVALID;
  wire [63:0] m_axi_rmem14___Stream2Mmap_14___mmap_ARADDR;
  wire [1:0] m_axi_rmem14___Stream2Mmap_14___mmap_ARBURST;
  wire [3:0] m_axi_rmem14___Stream2Mmap_14___mmap_ARCACHE;
  wire [0:0] m_axi_rmem14___Stream2Mmap_14___mmap_ARID;
  wire [7:0] m_axi_rmem14___Stream2Mmap_14___mmap_ARLEN;
  wire m_axi_rmem14___Stream2Mmap_14___mmap_ARLOCK;
  wire [2:0] m_axi_rmem14___Stream2Mmap_14___mmap_ARPROT;
  wire [3:0] m_axi_rmem14___Stream2Mmap_14___mmap_ARQOS;
  wire m_axi_rmem14___Stream2Mmap_14___mmap_ARREADY;
  wire [2:0] m_axi_rmem14___Stream2Mmap_14___mmap_ARSIZE;
  wire m_axi_rmem14___Stream2Mmap_14___mmap_ARVALID;
  wire [63:0] m_axi_rmem14___Stream2Mmap_14___mmap_AWADDR;
  wire [1:0] m_axi_rmem14___Stream2Mmap_14___mmap_AWBURST;
  wire [3:0] m_axi_rmem14___Stream2Mmap_14___mmap_AWCACHE;
  wire [0:0] m_axi_rmem14___Stream2Mmap_14___mmap_AWID;
  wire [7:0] m_axi_rmem14___Stream2Mmap_14___mmap_AWLEN;
  wire m_axi_rmem14___Stream2Mmap_14___mmap_AWLOCK;
  wire [2:0] m_axi_rmem14___Stream2Mmap_14___mmap_AWPROT;
  wire [3:0] m_axi_rmem14___Stream2Mmap_14___mmap_AWQOS;
  wire m_axi_rmem14___Stream2Mmap_14___mmap_AWREADY;
  wire [2:0] m_axi_rmem14___Stream2Mmap_14___mmap_AWSIZE;
  wire m_axi_rmem14___Stream2Mmap_14___mmap_AWVALID;
  wire [0:0] m_axi_rmem14___Stream2Mmap_14___mmap_BID;
  wire m_axi_rmem14___Stream2Mmap_14___mmap_BREADY;
  wire [1:0] m_axi_rmem14___Stream2Mmap_14___mmap_BRESP;
  wire m_axi_rmem14___Stream2Mmap_14___mmap_BVALID;
  wire [511:0] m_axi_rmem14___Stream2Mmap_14___mmap_RDATA;
  wire [0:0] m_axi_rmem14___Stream2Mmap_14___mmap_RID;
  wire m_axi_rmem14___Stream2Mmap_14___mmap_RLAST;
  wire m_axi_rmem14___Stream2Mmap_14___mmap_RREADY;
  wire [1:0] m_axi_rmem14___Stream2Mmap_14___mmap_RRESP;
  wire m_axi_rmem14___Stream2Mmap_14___mmap_RVALID;
  wire [511:0] m_axi_rmem14___Stream2Mmap_14___mmap_WDATA;
  wire m_axi_rmem14___Stream2Mmap_14___mmap_WLAST;
  wire m_axi_rmem14___Stream2Mmap_14___mmap_WREADY;
  wire [63:0] m_axi_rmem14___Stream2Mmap_14___mmap_WSTRB;
  wire m_axi_rmem14___Stream2Mmap_14___mmap_WVALID;
  wire [63:0] m_axi_rmem15___Mmap2Stream_15___mmap_ARADDR;
  wire [1:0] m_axi_rmem15___Mmap2Stream_15___mmap_ARBURST;
  wire [3:0] m_axi_rmem15___Mmap2Stream_15___mmap_ARCACHE;
  wire [0:0] m_axi_rmem15___Mmap2Stream_15___mmap_ARID;
  wire [7:0] m_axi_rmem15___Mmap2Stream_15___mmap_ARLEN;
  wire m_axi_rmem15___Mmap2Stream_15___mmap_ARLOCK;
  wire [2:0] m_axi_rmem15___Mmap2Stream_15___mmap_ARPROT;
  wire [3:0] m_axi_rmem15___Mmap2Stream_15___mmap_ARQOS;
  wire m_axi_rmem15___Mmap2Stream_15___mmap_ARREADY;
  wire [2:0] m_axi_rmem15___Mmap2Stream_15___mmap_ARSIZE;
  wire m_axi_rmem15___Mmap2Stream_15___mmap_ARVALID;
  wire [63:0] m_axi_rmem15___Mmap2Stream_15___mmap_AWADDR;
  wire [1:0] m_axi_rmem15___Mmap2Stream_15___mmap_AWBURST;
  wire [3:0] m_axi_rmem15___Mmap2Stream_15___mmap_AWCACHE;
  wire [0:0] m_axi_rmem15___Mmap2Stream_15___mmap_AWID;
  wire [7:0] m_axi_rmem15___Mmap2Stream_15___mmap_AWLEN;
  wire m_axi_rmem15___Mmap2Stream_15___mmap_AWLOCK;
  wire [2:0] m_axi_rmem15___Mmap2Stream_15___mmap_AWPROT;
  wire [3:0] m_axi_rmem15___Mmap2Stream_15___mmap_AWQOS;
  wire m_axi_rmem15___Mmap2Stream_15___mmap_AWREADY;
  wire [2:0] m_axi_rmem15___Mmap2Stream_15___mmap_AWSIZE;
  wire m_axi_rmem15___Mmap2Stream_15___mmap_AWVALID;
  wire [0:0] m_axi_rmem15___Mmap2Stream_15___mmap_BID;
  wire m_axi_rmem15___Mmap2Stream_15___mmap_BREADY;
  wire [1:0] m_axi_rmem15___Mmap2Stream_15___mmap_BRESP;
  wire m_axi_rmem15___Mmap2Stream_15___mmap_BVALID;
  wire [511:0] m_axi_rmem15___Mmap2Stream_15___mmap_RDATA;
  wire [0:0] m_axi_rmem15___Mmap2Stream_15___mmap_RID;
  wire m_axi_rmem15___Mmap2Stream_15___mmap_RLAST;
  wire m_axi_rmem15___Mmap2Stream_15___mmap_RREADY;
  wire [1:0] m_axi_rmem15___Mmap2Stream_15___mmap_RRESP;
  wire m_axi_rmem15___Mmap2Stream_15___mmap_RVALID;
  wire [511:0] m_axi_rmem15___Mmap2Stream_15___mmap_WDATA;
  wire m_axi_rmem15___Mmap2Stream_15___mmap_WLAST;
  wire m_axi_rmem15___Mmap2Stream_15___mmap_WREADY;
  wire [63:0] m_axi_rmem15___Mmap2Stream_15___mmap_WSTRB;
  wire m_axi_rmem15___Mmap2Stream_15___mmap_WVALID;
  wire [63:0] m_axi_rmem15___Stream2Mmap_15___mmap_ARADDR;
  wire [1:0] m_axi_rmem15___Stream2Mmap_15___mmap_ARBURST;
  wire [3:0] m_axi_rmem15___Stream2Mmap_15___mmap_ARCACHE;
  wire [0:0] m_axi_rmem15___Stream2Mmap_15___mmap_ARID;
  wire [7:0] m_axi_rmem15___Stream2Mmap_15___mmap_ARLEN;
  wire m_axi_rmem15___Stream2Mmap_15___mmap_ARLOCK;
  wire [2:0] m_axi_rmem15___Stream2Mmap_15___mmap_ARPROT;
  wire [3:0] m_axi_rmem15___Stream2Mmap_15___mmap_ARQOS;
  wire m_axi_rmem15___Stream2Mmap_15___mmap_ARREADY;
  wire [2:0] m_axi_rmem15___Stream2Mmap_15___mmap_ARSIZE;
  wire m_axi_rmem15___Stream2Mmap_15___mmap_ARVALID;
  wire [63:0] m_axi_rmem15___Stream2Mmap_15___mmap_AWADDR;
  wire [1:0] m_axi_rmem15___Stream2Mmap_15___mmap_AWBURST;
  wire [3:0] m_axi_rmem15___Stream2Mmap_15___mmap_AWCACHE;
  wire [0:0] m_axi_rmem15___Stream2Mmap_15___mmap_AWID;
  wire [7:0] m_axi_rmem15___Stream2Mmap_15___mmap_AWLEN;
  wire m_axi_rmem15___Stream2Mmap_15___mmap_AWLOCK;
  wire [2:0] m_axi_rmem15___Stream2Mmap_15___mmap_AWPROT;
  wire [3:0] m_axi_rmem15___Stream2Mmap_15___mmap_AWQOS;
  wire m_axi_rmem15___Stream2Mmap_15___mmap_AWREADY;
  wire [2:0] m_axi_rmem15___Stream2Mmap_15___mmap_AWSIZE;
  wire m_axi_rmem15___Stream2Mmap_15___mmap_AWVALID;
  wire [0:0] m_axi_rmem15___Stream2Mmap_15___mmap_BID;
  wire m_axi_rmem15___Stream2Mmap_15___mmap_BREADY;
  wire [1:0] m_axi_rmem15___Stream2Mmap_15___mmap_BRESP;
  wire m_axi_rmem15___Stream2Mmap_15___mmap_BVALID;
  wire [511:0] m_axi_rmem15___Stream2Mmap_15___mmap_RDATA;
  wire [0:0] m_axi_rmem15___Stream2Mmap_15___mmap_RID;
  wire m_axi_rmem15___Stream2Mmap_15___mmap_RLAST;
  wire m_axi_rmem15___Stream2Mmap_15___mmap_RREADY;
  wire [1:0] m_axi_rmem15___Stream2Mmap_15___mmap_RRESP;
  wire m_axi_rmem15___Stream2Mmap_15___mmap_RVALID;
  wire [511:0] m_axi_rmem15___Stream2Mmap_15___mmap_WDATA;
  wire m_axi_rmem15___Stream2Mmap_15___mmap_WLAST;
  wire m_axi_rmem15___Stream2Mmap_15___mmap_WREADY;
  wire [63:0] m_axi_rmem15___Stream2Mmap_15___mmap_WSTRB;
  wire m_axi_rmem15___Stream2Mmap_15___mmap_WVALID;
  wire [63:0] m_axi_rmem16___Mmap2Stream_16___mmap_ARADDR;
  wire [1:0] m_axi_rmem16___Mmap2Stream_16___mmap_ARBURST;
  wire [3:0] m_axi_rmem16___Mmap2Stream_16___mmap_ARCACHE;
  wire [0:0] m_axi_rmem16___Mmap2Stream_16___mmap_ARID;
  wire [7:0] m_axi_rmem16___Mmap2Stream_16___mmap_ARLEN;
  wire m_axi_rmem16___Mmap2Stream_16___mmap_ARLOCK;
  wire [2:0] m_axi_rmem16___Mmap2Stream_16___mmap_ARPROT;
  wire [3:0] m_axi_rmem16___Mmap2Stream_16___mmap_ARQOS;
  wire m_axi_rmem16___Mmap2Stream_16___mmap_ARREADY;
  wire [2:0] m_axi_rmem16___Mmap2Stream_16___mmap_ARSIZE;
  wire m_axi_rmem16___Mmap2Stream_16___mmap_ARVALID;
  wire [63:0] m_axi_rmem16___Mmap2Stream_16___mmap_AWADDR;
  wire [1:0] m_axi_rmem16___Mmap2Stream_16___mmap_AWBURST;
  wire [3:0] m_axi_rmem16___Mmap2Stream_16___mmap_AWCACHE;
  wire [0:0] m_axi_rmem16___Mmap2Stream_16___mmap_AWID;
  wire [7:0] m_axi_rmem16___Mmap2Stream_16___mmap_AWLEN;
  wire m_axi_rmem16___Mmap2Stream_16___mmap_AWLOCK;
  wire [2:0] m_axi_rmem16___Mmap2Stream_16___mmap_AWPROT;
  wire [3:0] m_axi_rmem16___Mmap2Stream_16___mmap_AWQOS;
  wire m_axi_rmem16___Mmap2Stream_16___mmap_AWREADY;
  wire [2:0] m_axi_rmem16___Mmap2Stream_16___mmap_AWSIZE;
  wire m_axi_rmem16___Mmap2Stream_16___mmap_AWVALID;
  wire [0:0] m_axi_rmem16___Mmap2Stream_16___mmap_BID;
  wire m_axi_rmem16___Mmap2Stream_16___mmap_BREADY;
  wire [1:0] m_axi_rmem16___Mmap2Stream_16___mmap_BRESP;
  wire m_axi_rmem16___Mmap2Stream_16___mmap_BVALID;
  wire [511:0] m_axi_rmem16___Mmap2Stream_16___mmap_RDATA;
  wire [0:0] m_axi_rmem16___Mmap2Stream_16___mmap_RID;
  wire m_axi_rmem16___Mmap2Stream_16___mmap_RLAST;
  wire m_axi_rmem16___Mmap2Stream_16___mmap_RREADY;
  wire [1:0] m_axi_rmem16___Mmap2Stream_16___mmap_RRESP;
  wire m_axi_rmem16___Mmap2Stream_16___mmap_RVALID;
  wire [511:0] m_axi_rmem16___Mmap2Stream_16___mmap_WDATA;
  wire m_axi_rmem16___Mmap2Stream_16___mmap_WLAST;
  wire m_axi_rmem16___Mmap2Stream_16___mmap_WREADY;
  wire [63:0] m_axi_rmem16___Mmap2Stream_16___mmap_WSTRB;
  wire m_axi_rmem16___Mmap2Stream_16___mmap_WVALID;
  wire [63:0] m_axi_rmem16___Stream2Mmap_16___mmap_ARADDR;
  wire [1:0] m_axi_rmem16___Stream2Mmap_16___mmap_ARBURST;
  wire [3:0] m_axi_rmem16___Stream2Mmap_16___mmap_ARCACHE;
  wire [0:0] m_axi_rmem16___Stream2Mmap_16___mmap_ARID;
  wire [7:0] m_axi_rmem16___Stream2Mmap_16___mmap_ARLEN;
  wire m_axi_rmem16___Stream2Mmap_16___mmap_ARLOCK;
  wire [2:0] m_axi_rmem16___Stream2Mmap_16___mmap_ARPROT;
  wire [3:0] m_axi_rmem16___Stream2Mmap_16___mmap_ARQOS;
  wire m_axi_rmem16___Stream2Mmap_16___mmap_ARREADY;
  wire [2:0] m_axi_rmem16___Stream2Mmap_16___mmap_ARSIZE;
  wire m_axi_rmem16___Stream2Mmap_16___mmap_ARVALID;
  wire [63:0] m_axi_rmem16___Stream2Mmap_16___mmap_AWADDR;
  wire [1:0] m_axi_rmem16___Stream2Mmap_16___mmap_AWBURST;
  wire [3:0] m_axi_rmem16___Stream2Mmap_16___mmap_AWCACHE;
  wire [0:0] m_axi_rmem16___Stream2Mmap_16___mmap_AWID;
  wire [7:0] m_axi_rmem16___Stream2Mmap_16___mmap_AWLEN;
  wire m_axi_rmem16___Stream2Mmap_16___mmap_AWLOCK;
  wire [2:0] m_axi_rmem16___Stream2Mmap_16___mmap_AWPROT;
  wire [3:0] m_axi_rmem16___Stream2Mmap_16___mmap_AWQOS;
  wire m_axi_rmem16___Stream2Mmap_16___mmap_AWREADY;
  wire [2:0] m_axi_rmem16___Stream2Mmap_16___mmap_AWSIZE;
  wire m_axi_rmem16___Stream2Mmap_16___mmap_AWVALID;
  wire [0:0] m_axi_rmem16___Stream2Mmap_16___mmap_BID;
  wire m_axi_rmem16___Stream2Mmap_16___mmap_BREADY;
  wire [1:0] m_axi_rmem16___Stream2Mmap_16___mmap_BRESP;
  wire m_axi_rmem16___Stream2Mmap_16___mmap_BVALID;
  wire [511:0] m_axi_rmem16___Stream2Mmap_16___mmap_RDATA;
  wire [0:0] m_axi_rmem16___Stream2Mmap_16___mmap_RID;
  wire m_axi_rmem16___Stream2Mmap_16___mmap_RLAST;
  wire m_axi_rmem16___Stream2Mmap_16___mmap_RREADY;
  wire [1:0] m_axi_rmem16___Stream2Mmap_16___mmap_RRESP;
  wire m_axi_rmem16___Stream2Mmap_16___mmap_RVALID;
  wire [511:0] m_axi_rmem16___Stream2Mmap_16___mmap_WDATA;
  wire m_axi_rmem16___Stream2Mmap_16___mmap_WLAST;
  wire m_axi_rmem16___Stream2Mmap_16___mmap_WREADY;
  wire [63:0] m_axi_rmem16___Stream2Mmap_16___mmap_WSTRB;
  wire m_axi_rmem16___Stream2Mmap_16___mmap_WVALID;
  wire [63:0] m_axi_rmem17___Mmap2Stream_17___mmap_ARADDR;
  wire [1:0] m_axi_rmem17___Mmap2Stream_17___mmap_ARBURST;
  wire [3:0] m_axi_rmem17___Mmap2Stream_17___mmap_ARCACHE;
  wire [0:0] m_axi_rmem17___Mmap2Stream_17___mmap_ARID;
  wire [7:0] m_axi_rmem17___Mmap2Stream_17___mmap_ARLEN;
  wire m_axi_rmem17___Mmap2Stream_17___mmap_ARLOCK;
  wire [2:0] m_axi_rmem17___Mmap2Stream_17___mmap_ARPROT;
  wire [3:0] m_axi_rmem17___Mmap2Stream_17___mmap_ARQOS;
  wire m_axi_rmem17___Mmap2Stream_17___mmap_ARREADY;
  wire [2:0] m_axi_rmem17___Mmap2Stream_17___mmap_ARSIZE;
  wire m_axi_rmem17___Mmap2Stream_17___mmap_ARVALID;
  wire [63:0] m_axi_rmem17___Mmap2Stream_17___mmap_AWADDR;
  wire [1:0] m_axi_rmem17___Mmap2Stream_17___mmap_AWBURST;
  wire [3:0] m_axi_rmem17___Mmap2Stream_17___mmap_AWCACHE;
  wire [0:0] m_axi_rmem17___Mmap2Stream_17___mmap_AWID;
  wire [7:0] m_axi_rmem17___Mmap2Stream_17___mmap_AWLEN;
  wire m_axi_rmem17___Mmap2Stream_17___mmap_AWLOCK;
  wire [2:0] m_axi_rmem17___Mmap2Stream_17___mmap_AWPROT;
  wire [3:0] m_axi_rmem17___Mmap2Stream_17___mmap_AWQOS;
  wire m_axi_rmem17___Mmap2Stream_17___mmap_AWREADY;
  wire [2:0] m_axi_rmem17___Mmap2Stream_17___mmap_AWSIZE;
  wire m_axi_rmem17___Mmap2Stream_17___mmap_AWVALID;
  wire [0:0] m_axi_rmem17___Mmap2Stream_17___mmap_BID;
  wire m_axi_rmem17___Mmap2Stream_17___mmap_BREADY;
  wire [1:0] m_axi_rmem17___Mmap2Stream_17___mmap_BRESP;
  wire m_axi_rmem17___Mmap2Stream_17___mmap_BVALID;
  wire [511:0] m_axi_rmem17___Mmap2Stream_17___mmap_RDATA;
  wire [0:0] m_axi_rmem17___Mmap2Stream_17___mmap_RID;
  wire m_axi_rmem17___Mmap2Stream_17___mmap_RLAST;
  wire m_axi_rmem17___Mmap2Stream_17___mmap_RREADY;
  wire [1:0] m_axi_rmem17___Mmap2Stream_17___mmap_RRESP;
  wire m_axi_rmem17___Mmap2Stream_17___mmap_RVALID;
  wire [511:0] m_axi_rmem17___Mmap2Stream_17___mmap_WDATA;
  wire m_axi_rmem17___Mmap2Stream_17___mmap_WLAST;
  wire m_axi_rmem17___Mmap2Stream_17___mmap_WREADY;
  wire [63:0] m_axi_rmem17___Mmap2Stream_17___mmap_WSTRB;
  wire m_axi_rmem17___Mmap2Stream_17___mmap_WVALID;
  wire [63:0] m_axi_rmem17___Stream2Mmap_17___mmap_ARADDR;
  wire [1:0] m_axi_rmem17___Stream2Mmap_17___mmap_ARBURST;
  wire [3:0] m_axi_rmem17___Stream2Mmap_17___mmap_ARCACHE;
  wire [0:0] m_axi_rmem17___Stream2Mmap_17___mmap_ARID;
  wire [7:0] m_axi_rmem17___Stream2Mmap_17___mmap_ARLEN;
  wire m_axi_rmem17___Stream2Mmap_17___mmap_ARLOCK;
  wire [2:0] m_axi_rmem17___Stream2Mmap_17___mmap_ARPROT;
  wire [3:0] m_axi_rmem17___Stream2Mmap_17___mmap_ARQOS;
  wire m_axi_rmem17___Stream2Mmap_17___mmap_ARREADY;
  wire [2:0] m_axi_rmem17___Stream2Mmap_17___mmap_ARSIZE;
  wire m_axi_rmem17___Stream2Mmap_17___mmap_ARVALID;
  wire [63:0] m_axi_rmem17___Stream2Mmap_17___mmap_AWADDR;
  wire [1:0] m_axi_rmem17___Stream2Mmap_17___mmap_AWBURST;
  wire [3:0] m_axi_rmem17___Stream2Mmap_17___mmap_AWCACHE;
  wire [0:0] m_axi_rmem17___Stream2Mmap_17___mmap_AWID;
  wire [7:0] m_axi_rmem17___Stream2Mmap_17___mmap_AWLEN;
  wire m_axi_rmem17___Stream2Mmap_17___mmap_AWLOCK;
  wire [2:0] m_axi_rmem17___Stream2Mmap_17___mmap_AWPROT;
  wire [3:0] m_axi_rmem17___Stream2Mmap_17___mmap_AWQOS;
  wire m_axi_rmem17___Stream2Mmap_17___mmap_AWREADY;
  wire [2:0] m_axi_rmem17___Stream2Mmap_17___mmap_AWSIZE;
  wire m_axi_rmem17___Stream2Mmap_17___mmap_AWVALID;
  wire [0:0] m_axi_rmem17___Stream2Mmap_17___mmap_BID;
  wire m_axi_rmem17___Stream2Mmap_17___mmap_BREADY;
  wire [1:0] m_axi_rmem17___Stream2Mmap_17___mmap_BRESP;
  wire m_axi_rmem17___Stream2Mmap_17___mmap_BVALID;
  wire [511:0] m_axi_rmem17___Stream2Mmap_17___mmap_RDATA;
  wire [0:0] m_axi_rmem17___Stream2Mmap_17___mmap_RID;
  wire m_axi_rmem17___Stream2Mmap_17___mmap_RLAST;
  wire m_axi_rmem17___Stream2Mmap_17___mmap_RREADY;
  wire [1:0] m_axi_rmem17___Stream2Mmap_17___mmap_RRESP;
  wire m_axi_rmem17___Stream2Mmap_17___mmap_RVALID;
  wire [511:0] m_axi_rmem17___Stream2Mmap_17___mmap_WDATA;
  wire m_axi_rmem17___Stream2Mmap_17___mmap_WLAST;
  wire m_axi_rmem17___Stream2Mmap_17___mmap_WREADY;
  wire [63:0] m_axi_rmem17___Stream2Mmap_17___mmap_WSTRB;
  wire m_axi_rmem17___Stream2Mmap_17___mmap_WVALID;
  wire [63:0] m_axi_rmem18___Mmap2Stream_18___mmap_ARADDR;
  wire [1:0] m_axi_rmem18___Mmap2Stream_18___mmap_ARBURST;
  wire [3:0] m_axi_rmem18___Mmap2Stream_18___mmap_ARCACHE;
  wire [0:0] m_axi_rmem18___Mmap2Stream_18___mmap_ARID;
  wire [7:0] m_axi_rmem18___Mmap2Stream_18___mmap_ARLEN;
  wire m_axi_rmem18___Mmap2Stream_18___mmap_ARLOCK;
  wire [2:0] m_axi_rmem18___Mmap2Stream_18___mmap_ARPROT;
  wire [3:0] m_axi_rmem18___Mmap2Stream_18___mmap_ARQOS;
  wire m_axi_rmem18___Mmap2Stream_18___mmap_ARREADY;
  wire [2:0] m_axi_rmem18___Mmap2Stream_18___mmap_ARSIZE;
  wire m_axi_rmem18___Mmap2Stream_18___mmap_ARVALID;
  wire [63:0] m_axi_rmem18___Mmap2Stream_18___mmap_AWADDR;
  wire [1:0] m_axi_rmem18___Mmap2Stream_18___mmap_AWBURST;
  wire [3:0] m_axi_rmem18___Mmap2Stream_18___mmap_AWCACHE;
  wire [0:0] m_axi_rmem18___Mmap2Stream_18___mmap_AWID;
  wire [7:0] m_axi_rmem18___Mmap2Stream_18___mmap_AWLEN;
  wire m_axi_rmem18___Mmap2Stream_18___mmap_AWLOCK;
  wire [2:0] m_axi_rmem18___Mmap2Stream_18___mmap_AWPROT;
  wire [3:0] m_axi_rmem18___Mmap2Stream_18___mmap_AWQOS;
  wire m_axi_rmem18___Mmap2Stream_18___mmap_AWREADY;
  wire [2:0] m_axi_rmem18___Mmap2Stream_18___mmap_AWSIZE;
  wire m_axi_rmem18___Mmap2Stream_18___mmap_AWVALID;
  wire [0:0] m_axi_rmem18___Mmap2Stream_18___mmap_BID;
  wire m_axi_rmem18___Mmap2Stream_18___mmap_BREADY;
  wire [1:0] m_axi_rmem18___Mmap2Stream_18___mmap_BRESP;
  wire m_axi_rmem18___Mmap2Stream_18___mmap_BVALID;
  wire [511:0] m_axi_rmem18___Mmap2Stream_18___mmap_RDATA;
  wire [0:0] m_axi_rmem18___Mmap2Stream_18___mmap_RID;
  wire m_axi_rmem18___Mmap2Stream_18___mmap_RLAST;
  wire m_axi_rmem18___Mmap2Stream_18___mmap_RREADY;
  wire [1:0] m_axi_rmem18___Mmap2Stream_18___mmap_RRESP;
  wire m_axi_rmem18___Mmap2Stream_18___mmap_RVALID;
  wire [511:0] m_axi_rmem18___Mmap2Stream_18___mmap_WDATA;
  wire m_axi_rmem18___Mmap2Stream_18___mmap_WLAST;
  wire m_axi_rmem18___Mmap2Stream_18___mmap_WREADY;
  wire [63:0] m_axi_rmem18___Mmap2Stream_18___mmap_WSTRB;
  wire m_axi_rmem18___Mmap2Stream_18___mmap_WVALID;
  wire [63:0] m_axi_rmem18___Stream2Mmap_18___mmap_ARADDR;
  wire [1:0] m_axi_rmem18___Stream2Mmap_18___mmap_ARBURST;
  wire [3:0] m_axi_rmem18___Stream2Mmap_18___mmap_ARCACHE;
  wire [0:0] m_axi_rmem18___Stream2Mmap_18___mmap_ARID;
  wire [7:0] m_axi_rmem18___Stream2Mmap_18___mmap_ARLEN;
  wire m_axi_rmem18___Stream2Mmap_18___mmap_ARLOCK;
  wire [2:0] m_axi_rmem18___Stream2Mmap_18___mmap_ARPROT;
  wire [3:0] m_axi_rmem18___Stream2Mmap_18___mmap_ARQOS;
  wire m_axi_rmem18___Stream2Mmap_18___mmap_ARREADY;
  wire [2:0] m_axi_rmem18___Stream2Mmap_18___mmap_ARSIZE;
  wire m_axi_rmem18___Stream2Mmap_18___mmap_ARVALID;
  wire [63:0] m_axi_rmem18___Stream2Mmap_18___mmap_AWADDR;
  wire [1:0] m_axi_rmem18___Stream2Mmap_18___mmap_AWBURST;
  wire [3:0] m_axi_rmem18___Stream2Mmap_18___mmap_AWCACHE;
  wire [0:0] m_axi_rmem18___Stream2Mmap_18___mmap_AWID;
  wire [7:0] m_axi_rmem18___Stream2Mmap_18___mmap_AWLEN;
  wire m_axi_rmem18___Stream2Mmap_18___mmap_AWLOCK;
  wire [2:0] m_axi_rmem18___Stream2Mmap_18___mmap_AWPROT;
  wire [3:0] m_axi_rmem18___Stream2Mmap_18___mmap_AWQOS;
  wire m_axi_rmem18___Stream2Mmap_18___mmap_AWREADY;
  wire [2:0] m_axi_rmem18___Stream2Mmap_18___mmap_AWSIZE;
  wire m_axi_rmem18___Stream2Mmap_18___mmap_AWVALID;
  wire [0:0] m_axi_rmem18___Stream2Mmap_18___mmap_BID;
  wire m_axi_rmem18___Stream2Mmap_18___mmap_BREADY;
  wire [1:0] m_axi_rmem18___Stream2Mmap_18___mmap_BRESP;
  wire m_axi_rmem18___Stream2Mmap_18___mmap_BVALID;
  wire [511:0] m_axi_rmem18___Stream2Mmap_18___mmap_RDATA;
  wire [0:0] m_axi_rmem18___Stream2Mmap_18___mmap_RID;
  wire m_axi_rmem18___Stream2Mmap_18___mmap_RLAST;
  wire m_axi_rmem18___Stream2Mmap_18___mmap_RREADY;
  wire [1:0] m_axi_rmem18___Stream2Mmap_18___mmap_RRESP;
  wire m_axi_rmem18___Stream2Mmap_18___mmap_RVALID;
  wire [511:0] m_axi_rmem18___Stream2Mmap_18___mmap_WDATA;
  wire m_axi_rmem18___Stream2Mmap_18___mmap_WLAST;
  wire m_axi_rmem18___Stream2Mmap_18___mmap_WREADY;
  wire [63:0] m_axi_rmem18___Stream2Mmap_18___mmap_WSTRB;
  wire m_axi_rmem18___Stream2Mmap_18___mmap_WVALID;
  wire [63:0] m_axi_rmem19___Mmap2Stream_19___mmap_ARADDR;
  wire [1:0] m_axi_rmem19___Mmap2Stream_19___mmap_ARBURST;
  wire [3:0] m_axi_rmem19___Mmap2Stream_19___mmap_ARCACHE;
  wire [0:0] m_axi_rmem19___Mmap2Stream_19___mmap_ARID;
  wire [7:0] m_axi_rmem19___Mmap2Stream_19___mmap_ARLEN;
  wire m_axi_rmem19___Mmap2Stream_19___mmap_ARLOCK;
  wire [2:0] m_axi_rmem19___Mmap2Stream_19___mmap_ARPROT;
  wire [3:0] m_axi_rmem19___Mmap2Stream_19___mmap_ARQOS;
  wire m_axi_rmem19___Mmap2Stream_19___mmap_ARREADY;
  wire [2:0] m_axi_rmem19___Mmap2Stream_19___mmap_ARSIZE;
  wire m_axi_rmem19___Mmap2Stream_19___mmap_ARVALID;
  wire [63:0] m_axi_rmem19___Mmap2Stream_19___mmap_AWADDR;
  wire [1:0] m_axi_rmem19___Mmap2Stream_19___mmap_AWBURST;
  wire [3:0] m_axi_rmem19___Mmap2Stream_19___mmap_AWCACHE;
  wire [0:0] m_axi_rmem19___Mmap2Stream_19___mmap_AWID;
  wire [7:0] m_axi_rmem19___Mmap2Stream_19___mmap_AWLEN;
  wire m_axi_rmem19___Mmap2Stream_19___mmap_AWLOCK;
  wire [2:0] m_axi_rmem19___Mmap2Stream_19___mmap_AWPROT;
  wire [3:0] m_axi_rmem19___Mmap2Stream_19___mmap_AWQOS;
  wire m_axi_rmem19___Mmap2Stream_19___mmap_AWREADY;
  wire [2:0] m_axi_rmem19___Mmap2Stream_19___mmap_AWSIZE;
  wire m_axi_rmem19___Mmap2Stream_19___mmap_AWVALID;
  wire [0:0] m_axi_rmem19___Mmap2Stream_19___mmap_BID;
  wire m_axi_rmem19___Mmap2Stream_19___mmap_BREADY;
  wire [1:0] m_axi_rmem19___Mmap2Stream_19___mmap_BRESP;
  wire m_axi_rmem19___Mmap2Stream_19___mmap_BVALID;
  wire [511:0] m_axi_rmem19___Mmap2Stream_19___mmap_RDATA;
  wire [0:0] m_axi_rmem19___Mmap2Stream_19___mmap_RID;
  wire m_axi_rmem19___Mmap2Stream_19___mmap_RLAST;
  wire m_axi_rmem19___Mmap2Stream_19___mmap_RREADY;
  wire [1:0] m_axi_rmem19___Mmap2Stream_19___mmap_RRESP;
  wire m_axi_rmem19___Mmap2Stream_19___mmap_RVALID;
  wire [511:0] m_axi_rmem19___Mmap2Stream_19___mmap_WDATA;
  wire m_axi_rmem19___Mmap2Stream_19___mmap_WLAST;
  wire m_axi_rmem19___Mmap2Stream_19___mmap_WREADY;
  wire [63:0] m_axi_rmem19___Mmap2Stream_19___mmap_WSTRB;
  wire m_axi_rmem19___Mmap2Stream_19___mmap_WVALID;
  wire [63:0] m_axi_rmem19___Stream2Mmap_19___mmap_ARADDR;
  wire [1:0] m_axi_rmem19___Stream2Mmap_19___mmap_ARBURST;
  wire [3:0] m_axi_rmem19___Stream2Mmap_19___mmap_ARCACHE;
  wire [0:0] m_axi_rmem19___Stream2Mmap_19___mmap_ARID;
  wire [7:0] m_axi_rmem19___Stream2Mmap_19___mmap_ARLEN;
  wire m_axi_rmem19___Stream2Mmap_19___mmap_ARLOCK;
  wire [2:0] m_axi_rmem19___Stream2Mmap_19___mmap_ARPROT;
  wire [3:0] m_axi_rmem19___Stream2Mmap_19___mmap_ARQOS;
  wire m_axi_rmem19___Stream2Mmap_19___mmap_ARREADY;
  wire [2:0] m_axi_rmem19___Stream2Mmap_19___mmap_ARSIZE;
  wire m_axi_rmem19___Stream2Mmap_19___mmap_ARVALID;
  wire [63:0] m_axi_rmem19___Stream2Mmap_19___mmap_AWADDR;
  wire [1:0] m_axi_rmem19___Stream2Mmap_19___mmap_AWBURST;
  wire [3:0] m_axi_rmem19___Stream2Mmap_19___mmap_AWCACHE;
  wire [0:0] m_axi_rmem19___Stream2Mmap_19___mmap_AWID;
  wire [7:0] m_axi_rmem19___Stream2Mmap_19___mmap_AWLEN;
  wire m_axi_rmem19___Stream2Mmap_19___mmap_AWLOCK;
  wire [2:0] m_axi_rmem19___Stream2Mmap_19___mmap_AWPROT;
  wire [3:0] m_axi_rmem19___Stream2Mmap_19___mmap_AWQOS;
  wire m_axi_rmem19___Stream2Mmap_19___mmap_AWREADY;
  wire [2:0] m_axi_rmem19___Stream2Mmap_19___mmap_AWSIZE;
  wire m_axi_rmem19___Stream2Mmap_19___mmap_AWVALID;
  wire [0:0] m_axi_rmem19___Stream2Mmap_19___mmap_BID;
  wire m_axi_rmem19___Stream2Mmap_19___mmap_BREADY;
  wire [1:0] m_axi_rmem19___Stream2Mmap_19___mmap_BRESP;
  wire m_axi_rmem19___Stream2Mmap_19___mmap_BVALID;
  wire [511:0] m_axi_rmem19___Stream2Mmap_19___mmap_RDATA;
  wire [0:0] m_axi_rmem19___Stream2Mmap_19___mmap_RID;
  wire m_axi_rmem19___Stream2Mmap_19___mmap_RLAST;
  wire m_axi_rmem19___Stream2Mmap_19___mmap_RREADY;
  wire [1:0] m_axi_rmem19___Stream2Mmap_19___mmap_RRESP;
  wire m_axi_rmem19___Stream2Mmap_19___mmap_RVALID;
  wire [511:0] m_axi_rmem19___Stream2Mmap_19___mmap_WDATA;
  wire m_axi_rmem19___Stream2Mmap_19___mmap_WLAST;
  wire m_axi_rmem19___Stream2Mmap_19___mmap_WREADY;
  wire [63:0] m_axi_rmem19___Stream2Mmap_19___mmap_WSTRB;
  wire m_axi_rmem19___Stream2Mmap_19___mmap_WVALID;
  wire [63:0] m_axi_rmem20___Mmap2Stream_20___mmap_ARADDR;
  wire [1:0] m_axi_rmem20___Mmap2Stream_20___mmap_ARBURST;
  wire [3:0] m_axi_rmem20___Mmap2Stream_20___mmap_ARCACHE;
  wire [0:0] m_axi_rmem20___Mmap2Stream_20___mmap_ARID;
  wire [7:0] m_axi_rmem20___Mmap2Stream_20___mmap_ARLEN;
  wire m_axi_rmem20___Mmap2Stream_20___mmap_ARLOCK;
  wire [2:0] m_axi_rmem20___Mmap2Stream_20___mmap_ARPROT;
  wire [3:0] m_axi_rmem20___Mmap2Stream_20___mmap_ARQOS;
  wire m_axi_rmem20___Mmap2Stream_20___mmap_ARREADY;
  wire [2:0] m_axi_rmem20___Mmap2Stream_20___mmap_ARSIZE;
  wire m_axi_rmem20___Mmap2Stream_20___mmap_ARVALID;
  wire [63:0] m_axi_rmem20___Mmap2Stream_20___mmap_AWADDR;
  wire [1:0] m_axi_rmem20___Mmap2Stream_20___mmap_AWBURST;
  wire [3:0] m_axi_rmem20___Mmap2Stream_20___mmap_AWCACHE;
  wire [0:0] m_axi_rmem20___Mmap2Stream_20___mmap_AWID;
  wire [7:0] m_axi_rmem20___Mmap2Stream_20___mmap_AWLEN;
  wire m_axi_rmem20___Mmap2Stream_20___mmap_AWLOCK;
  wire [2:0] m_axi_rmem20___Mmap2Stream_20___mmap_AWPROT;
  wire [3:0] m_axi_rmem20___Mmap2Stream_20___mmap_AWQOS;
  wire m_axi_rmem20___Mmap2Stream_20___mmap_AWREADY;
  wire [2:0] m_axi_rmem20___Mmap2Stream_20___mmap_AWSIZE;
  wire m_axi_rmem20___Mmap2Stream_20___mmap_AWVALID;
  wire [0:0] m_axi_rmem20___Mmap2Stream_20___mmap_BID;
  wire m_axi_rmem20___Mmap2Stream_20___mmap_BREADY;
  wire [1:0] m_axi_rmem20___Mmap2Stream_20___mmap_BRESP;
  wire m_axi_rmem20___Mmap2Stream_20___mmap_BVALID;
  wire [511:0] m_axi_rmem20___Mmap2Stream_20___mmap_RDATA;
  wire [0:0] m_axi_rmem20___Mmap2Stream_20___mmap_RID;
  wire m_axi_rmem20___Mmap2Stream_20___mmap_RLAST;
  wire m_axi_rmem20___Mmap2Stream_20___mmap_RREADY;
  wire [1:0] m_axi_rmem20___Mmap2Stream_20___mmap_RRESP;
  wire m_axi_rmem20___Mmap2Stream_20___mmap_RVALID;
  wire [511:0] m_axi_rmem20___Mmap2Stream_20___mmap_WDATA;
  wire m_axi_rmem20___Mmap2Stream_20___mmap_WLAST;
  wire m_axi_rmem20___Mmap2Stream_20___mmap_WREADY;
  wire [63:0] m_axi_rmem20___Mmap2Stream_20___mmap_WSTRB;
  wire m_axi_rmem20___Mmap2Stream_20___mmap_WVALID;
  wire [63:0] m_axi_rmem20___Stream2Mmap_20___mmap_ARADDR;
  wire [1:0] m_axi_rmem20___Stream2Mmap_20___mmap_ARBURST;
  wire [3:0] m_axi_rmem20___Stream2Mmap_20___mmap_ARCACHE;
  wire [0:0] m_axi_rmem20___Stream2Mmap_20___mmap_ARID;
  wire [7:0] m_axi_rmem20___Stream2Mmap_20___mmap_ARLEN;
  wire m_axi_rmem20___Stream2Mmap_20___mmap_ARLOCK;
  wire [2:0] m_axi_rmem20___Stream2Mmap_20___mmap_ARPROT;
  wire [3:0] m_axi_rmem20___Stream2Mmap_20___mmap_ARQOS;
  wire m_axi_rmem20___Stream2Mmap_20___mmap_ARREADY;
  wire [2:0] m_axi_rmem20___Stream2Mmap_20___mmap_ARSIZE;
  wire m_axi_rmem20___Stream2Mmap_20___mmap_ARVALID;
  wire [63:0] m_axi_rmem20___Stream2Mmap_20___mmap_AWADDR;
  wire [1:0] m_axi_rmem20___Stream2Mmap_20___mmap_AWBURST;
  wire [3:0] m_axi_rmem20___Stream2Mmap_20___mmap_AWCACHE;
  wire [0:0] m_axi_rmem20___Stream2Mmap_20___mmap_AWID;
  wire [7:0] m_axi_rmem20___Stream2Mmap_20___mmap_AWLEN;
  wire m_axi_rmem20___Stream2Mmap_20___mmap_AWLOCK;
  wire [2:0] m_axi_rmem20___Stream2Mmap_20___mmap_AWPROT;
  wire [3:0] m_axi_rmem20___Stream2Mmap_20___mmap_AWQOS;
  wire m_axi_rmem20___Stream2Mmap_20___mmap_AWREADY;
  wire [2:0] m_axi_rmem20___Stream2Mmap_20___mmap_AWSIZE;
  wire m_axi_rmem20___Stream2Mmap_20___mmap_AWVALID;
  wire [0:0] m_axi_rmem20___Stream2Mmap_20___mmap_BID;
  wire m_axi_rmem20___Stream2Mmap_20___mmap_BREADY;
  wire [1:0] m_axi_rmem20___Stream2Mmap_20___mmap_BRESP;
  wire m_axi_rmem20___Stream2Mmap_20___mmap_BVALID;
  wire [511:0] m_axi_rmem20___Stream2Mmap_20___mmap_RDATA;
  wire [0:0] m_axi_rmem20___Stream2Mmap_20___mmap_RID;
  wire m_axi_rmem20___Stream2Mmap_20___mmap_RLAST;
  wire m_axi_rmem20___Stream2Mmap_20___mmap_RREADY;
  wire [1:0] m_axi_rmem20___Stream2Mmap_20___mmap_RRESP;
  wire m_axi_rmem20___Stream2Mmap_20___mmap_RVALID;
  wire [511:0] m_axi_rmem20___Stream2Mmap_20___mmap_WDATA;
  wire m_axi_rmem20___Stream2Mmap_20___mmap_WLAST;
  wire m_axi_rmem20___Stream2Mmap_20___mmap_WREADY;
  wire [63:0] m_axi_rmem20___Stream2Mmap_20___mmap_WSTRB;
  wire m_axi_rmem20___Stream2Mmap_20___mmap_WVALID;
  wire [63:0] m_axi_rmem21___Mmap2Stream_21___mmap_ARADDR;
  wire [1:0] m_axi_rmem21___Mmap2Stream_21___mmap_ARBURST;
  wire [3:0] m_axi_rmem21___Mmap2Stream_21___mmap_ARCACHE;
  wire [0:0] m_axi_rmem21___Mmap2Stream_21___mmap_ARID;
  wire [7:0] m_axi_rmem21___Mmap2Stream_21___mmap_ARLEN;
  wire m_axi_rmem21___Mmap2Stream_21___mmap_ARLOCK;
  wire [2:0] m_axi_rmem21___Mmap2Stream_21___mmap_ARPROT;
  wire [3:0] m_axi_rmem21___Mmap2Stream_21___mmap_ARQOS;
  wire m_axi_rmem21___Mmap2Stream_21___mmap_ARREADY;
  wire [2:0] m_axi_rmem21___Mmap2Stream_21___mmap_ARSIZE;
  wire m_axi_rmem21___Mmap2Stream_21___mmap_ARVALID;
  wire [63:0] m_axi_rmem21___Mmap2Stream_21___mmap_AWADDR;
  wire [1:0] m_axi_rmem21___Mmap2Stream_21___mmap_AWBURST;
  wire [3:0] m_axi_rmem21___Mmap2Stream_21___mmap_AWCACHE;
  wire [0:0] m_axi_rmem21___Mmap2Stream_21___mmap_AWID;
  wire [7:0] m_axi_rmem21___Mmap2Stream_21___mmap_AWLEN;
  wire m_axi_rmem21___Mmap2Stream_21___mmap_AWLOCK;
  wire [2:0] m_axi_rmem21___Mmap2Stream_21___mmap_AWPROT;
  wire [3:0] m_axi_rmem21___Mmap2Stream_21___mmap_AWQOS;
  wire m_axi_rmem21___Mmap2Stream_21___mmap_AWREADY;
  wire [2:0] m_axi_rmem21___Mmap2Stream_21___mmap_AWSIZE;
  wire m_axi_rmem21___Mmap2Stream_21___mmap_AWVALID;
  wire [0:0] m_axi_rmem21___Mmap2Stream_21___mmap_BID;
  wire m_axi_rmem21___Mmap2Stream_21___mmap_BREADY;
  wire [1:0] m_axi_rmem21___Mmap2Stream_21___mmap_BRESP;
  wire m_axi_rmem21___Mmap2Stream_21___mmap_BVALID;
  wire [511:0] m_axi_rmem21___Mmap2Stream_21___mmap_RDATA;
  wire [0:0] m_axi_rmem21___Mmap2Stream_21___mmap_RID;
  wire m_axi_rmem21___Mmap2Stream_21___mmap_RLAST;
  wire m_axi_rmem21___Mmap2Stream_21___mmap_RREADY;
  wire [1:0] m_axi_rmem21___Mmap2Stream_21___mmap_RRESP;
  wire m_axi_rmem21___Mmap2Stream_21___mmap_RVALID;
  wire [511:0] m_axi_rmem21___Mmap2Stream_21___mmap_WDATA;
  wire m_axi_rmem21___Mmap2Stream_21___mmap_WLAST;
  wire m_axi_rmem21___Mmap2Stream_21___mmap_WREADY;
  wire [63:0] m_axi_rmem21___Mmap2Stream_21___mmap_WSTRB;
  wire m_axi_rmem21___Mmap2Stream_21___mmap_WVALID;
  wire [63:0] m_axi_rmem21___Stream2Mmap_21___mmap_ARADDR;
  wire [1:0] m_axi_rmem21___Stream2Mmap_21___mmap_ARBURST;
  wire [3:0] m_axi_rmem21___Stream2Mmap_21___mmap_ARCACHE;
  wire [0:0] m_axi_rmem21___Stream2Mmap_21___mmap_ARID;
  wire [7:0] m_axi_rmem21___Stream2Mmap_21___mmap_ARLEN;
  wire m_axi_rmem21___Stream2Mmap_21___mmap_ARLOCK;
  wire [2:0] m_axi_rmem21___Stream2Mmap_21___mmap_ARPROT;
  wire [3:0] m_axi_rmem21___Stream2Mmap_21___mmap_ARQOS;
  wire m_axi_rmem21___Stream2Mmap_21___mmap_ARREADY;
  wire [2:0] m_axi_rmem21___Stream2Mmap_21___mmap_ARSIZE;
  wire m_axi_rmem21___Stream2Mmap_21___mmap_ARVALID;
  wire [63:0] m_axi_rmem21___Stream2Mmap_21___mmap_AWADDR;
  wire [1:0] m_axi_rmem21___Stream2Mmap_21___mmap_AWBURST;
  wire [3:0] m_axi_rmem21___Stream2Mmap_21___mmap_AWCACHE;
  wire [0:0] m_axi_rmem21___Stream2Mmap_21___mmap_AWID;
  wire [7:0] m_axi_rmem21___Stream2Mmap_21___mmap_AWLEN;
  wire m_axi_rmem21___Stream2Mmap_21___mmap_AWLOCK;
  wire [2:0] m_axi_rmem21___Stream2Mmap_21___mmap_AWPROT;
  wire [3:0] m_axi_rmem21___Stream2Mmap_21___mmap_AWQOS;
  wire m_axi_rmem21___Stream2Mmap_21___mmap_AWREADY;
  wire [2:0] m_axi_rmem21___Stream2Mmap_21___mmap_AWSIZE;
  wire m_axi_rmem21___Stream2Mmap_21___mmap_AWVALID;
  wire [0:0] m_axi_rmem21___Stream2Mmap_21___mmap_BID;
  wire m_axi_rmem21___Stream2Mmap_21___mmap_BREADY;
  wire [1:0] m_axi_rmem21___Stream2Mmap_21___mmap_BRESP;
  wire m_axi_rmem21___Stream2Mmap_21___mmap_BVALID;
  wire [511:0] m_axi_rmem21___Stream2Mmap_21___mmap_RDATA;
  wire [0:0] m_axi_rmem21___Stream2Mmap_21___mmap_RID;
  wire m_axi_rmem21___Stream2Mmap_21___mmap_RLAST;
  wire m_axi_rmem21___Stream2Mmap_21___mmap_RREADY;
  wire [1:0] m_axi_rmem21___Stream2Mmap_21___mmap_RRESP;
  wire m_axi_rmem21___Stream2Mmap_21___mmap_RVALID;
  wire [511:0] m_axi_rmem21___Stream2Mmap_21___mmap_WDATA;
  wire m_axi_rmem21___Stream2Mmap_21___mmap_WLAST;
  wire m_axi_rmem21___Stream2Mmap_21___mmap_WREADY;
  wire [63:0] m_axi_rmem21___Stream2Mmap_21___mmap_WSTRB;
  wire m_axi_rmem21___Stream2Mmap_21___mmap_WVALID;
  wire [63:0] m_axi_rmem22___Mmap2Stream_22___mmap_ARADDR;
  wire [1:0] m_axi_rmem22___Mmap2Stream_22___mmap_ARBURST;
  wire [3:0] m_axi_rmem22___Mmap2Stream_22___mmap_ARCACHE;
  wire [0:0] m_axi_rmem22___Mmap2Stream_22___mmap_ARID;
  wire [7:0] m_axi_rmem22___Mmap2Stream_22___mmap_ARLEN;
  wire m_axi_rmem22___Mmap2Stream_22___mmap_ARLOCK;
  wire [2:0] m_axi_rmem22___Mmap2Stream_22___mmap_ARPROT;
  wire [3:0] m_axi_rmem22___Mmap2Stream_22___mmap_ARQOS;
  wire m_axi_rmem22___Mmap2Stream_22___mmap_ARREADY;
  wire [2:0] m_axi_rmem22___Mmap2Stream_22___mmap_ARSIZE;
  wire m_axi_rmem22___Mmap2Stream_22___mmap_ARVALID;
  wire [63:0] m_axi_rmem22___Mmap2Stream_22___mmap_AWADDR;
  wire [1:0] m_axi_rmem22___Mmap2Stream_22___mmap_AWBURST;
  wire [3:0] m_axi_rmem22___Mmap2Stream_22___mmap_AWCACHE;
  wire [0:0] m_axi_rmem22___Mmap2Stream_22___mmap_AWID;
  wire [7:0] m_axi_rmem22___Mmap2Stream_22___mmap_AWLEN;
  wire m_axi_rmem22___Mmap2Stream_22___mmap_AWLOCK;
  wire [2:0] m_axi_rmem22___Mmap2Stream_22___mmap_AWPROT;
  wire [3:0] m_axi_rmem22___Mmap2Stream_22___mmap_AWQOS;
  wire m_axi_rmem22___Mmap2Stream_22___mmap_AWREADY;
  wire [2:0] m_axi_rmem22___Mmap2Stream_22___mmap_AWSIZE;
  wire m_axi_rmem22___Mmap2Stream_22___mmap_AWVALID;
  wire [0:0] m_axi_rmem22___Mmap2Stream_22___mmap_BID;
  wire m_axi_rmem22___Mmap2Stream_22___mmap_BREADY;
  wire [1:0] m_axi_rmem22___Mmap2Stream_22___mmap_BRESP;
  wire m_axi_rmem22___Mmap2Stream_22___mmap_BVALID;
  wire [511:0] m_axi_rmem22___Mmap2Stream_22___mmap_RDATA;
  wire [0:0] m_axi_rmem22___Mmap2Stream_22___mmap_RID;
  wire m_axi_rmem22___Mmap2Stream_22___mmap_RLAST;
  wire m_axi_rmem22___Mmap2Stream_22___mmap_RREADY;
  wire [1:0] m_axi_rmem22___Mmap2Stream_22___mmap_RRESP;
  wire m_axi_rmem22___Mmap2Stream_22___mmap_RVALID;
  wire [511:0] m_axi_rmem22___Mmap2Stream_22___mmap_WDATA;
  wire m_axi_rmem22___Mmap2Stream_22___mmap_WLAST;
  wire m_axi_rmem22___Mmap2Stream_22___mmap_WREADY;
  wire [63:0] m_axi_rmem22___Mmap2Stream_22___mmap_WSTRB;
  wire m_axi_rmem22___Mmap2Stream_22___mmap_WVALID;
  wire [63:0] m_axi_rmem22___Stream2Mmap_22___mmap_ARADDR;
  wire [1:0] m_axi_rmem22___Stream2Mmap_22___mmap_ARBURST;
  wire [3:0] m_axi_rmem22___Stream2Mmap_22___mmap_ARCACHE;
  wire [0:0] m_axi_rmem22___Stream2Mmap_22___mmap_ARID;
  wire [7:0] m_axi_rmem22___Stream2Mmap_22___mmap_ARLEN;
  wire m_axi_rmem22___Stream2Mmap_22___mmap_ARLOCK;
  wire [2:0] m_axi_rmem22___Stream2Mmap_22___mmap_ARPROT;
  wire [3:0] m_axi_rmem22___Stream2Mmap_22___mmap_ARQOS;
  wire m_axi_rmem22___Stream2Mmap_22___mmap_ARREADY;
  wire [2:0] m_axi_rmem22___Stream2Mmap_22___mmap_ARSIZE;
  wire m_axi_rmem22___Stream2Mmap_22___mmap_ARVALID;
  wire [63:0] m_axi_rmem22___Stream2Mmap_22___mmap_AWADDR;
  wire [1:0] m_axi_rmem22___Stream2Mmap_22___mmap_AWBURST;
  wire [3:0] m_axi_rmem22___Stream2Mmap_22___mmap_AWCACHE;
  wire [0:0] m_axi_rmem22___Stream2Mmap_22___mmap_AWID;
  wire [7:0] m_axi_rmem22___Stream2Mmap_22___mmap_AWLEN;
  wire m_axi_rmem22___Stream2Mmap_22___mmap_AWLOCK;
  wire [2:0] m_axi_rmem22___Stream2Mmap_22___mmap_AWPROT;
  wire [3:0] m_axi_rmem22___Stream2Mmap_22___mmap_AWQOS;
  wire m_axi_rmem22___Stream2Mmap_22___mmap_AWREADY;
  wire [2:0] m_axi_rmem22___Stream2Mmap_22___mmap_AWSIZE;
  wire m_axi_rmem22___Stream2Mmap_22___mmap_AWVALID;
  wire [0:0] m_axi_rmem22___Stream2Mmap_22___mmap_BID;
  wire m_axi_rmem22___Stream2Mmap_22___mmap_BREADY;
  wire [1:0] m_axi_rmem22___Stream2Mmap_22___mmap_BRESP;
  wire m_axi_rmem22___Stream2Mmap_22___mmap_BVALID;
  wire [511:0] m_axi_rmem22___Stream2Mmap_22___mmap_RDATA;
  wire [0:0] m_axi_rmem22___Stream2Mmap_22___mmap_RID;
  wire m_axi_rmem22___Stream2Mmap_22___mmap_RLAST;
  wire m_axi_rmem22___Stream2Mmap_22___mmap_RREADY;
  wire [1:0] m_axi_rmem22___Stream2Mmap_22___mmap_RRESP;
  wire m_axi_rmem22___Stream2Mmap_22___mmap_RVALID;
  wire [511:0] m_axi_rmem22___Stream2Mmap_22___mmap_WDATA;
  wire m_axi_rmem22___Stream2Mmap_22___mmap_WLAST;
  wire m_axi_rmem22___Stream2Mmap_22___mmap_WREADY;
  wire [63:0] m_axi_rmem22___Stream2Mmap_22___mmap_WSTRB;
  wire m_axi_rmem22___Stream2Mmap_22___mmap_WVALID;
  wire [63:0] m_axi_rmem23___Mmap2Stream_23___mmap_ARADDR;
  wire [1:0] m_axi_rmem23___Mmap2Stream_23___mmap_ARBURST;
  wire [3:0] m_axi_rmem23___Mmap2Stream_23___mmap_ARCACHE;
  wire [0:0] m_axi_rmem23___Mmap2Stream_23___mmap_ARID;
  wire [7:0] m_axi_rmem23___Mmap2Stream_23___mmap_ARLEN;
  wire m_axi_rmem23___Mmap2Stream_23___mmap_ARLOCK;
  wire [2:0] m_axi_rmem23___Mmap2Stream_23___mmap_ARPROT;
  wire [3:0] m_axi_rmem23___Mmap2Stream_23___mmap_ARQOS;
  wire m_axi_rmem23___Mmap2Stream_23___mmap_ARREADY;
  wire [2:0] m_axi_rmem23___Mmap2Stream_23___mmap_ARSIZE;
  wire m_axi_rmem23___Mmap2Stream_23___mmap_ARVALID;
  wire [63:0] m_axi_rmem23___Mmap2Stream_23___mmap_AWADDR;
  wire [1:0] m_axi_rmem23___Mmap2Stream_23___mmap_AWBURST;
  wire [3:0] m_axi_rmem23___Mmap2Stream_23___mmap_AWCACHE;
  wire [0:0] m_axi_rmem23___Mmap2Stream_23___mmap_AWID;
  wire [7:0] m_axi_rmem23___Mmap2Stream_23___mmap_AWLEN;
  wire m_axi_rmem23___Mmap2Stream_23___mmap_AWLOCK;
  wire [2:0] m_axi_rmem23___Mmap2Stream_23___mmap_AWPROT;
  wire [3:0] m_axi_rmem23___Mmap2Stream_23___mmap_AWQOS;
  wire m_axi_rmem23___Mmap2Stream_23___mmap_AWREADY;
  wire [2:0] m_axi_rmem23___Mmap2Stream_23___mmap_AWSIZE;
  wire m_axi_rmem23___Mmap2Stream_23___mmap_AWVALID;
  wire [0:0] m_axi_rmem23___Mmap2Stream_23___mmap_BID;
  wire m_axi_rmem23___Mmap2Stream_23___mmap_BREADY;
  wire [1:0] m_axi_rmem23___Mmap2Stream_23___mmap_BRESP;
  wire m_axi_rmem23___Mmap2Stream_23___mmap_BVALID;
  wire [511:0] m_axi_rmem23___Mmap2Stream_23___mmap_RDATA;
  wire [0:0] m_axi_rmem23___Mmap2Stream_23___mmap_RID;
  wire m_axi_rmem23___Mmap2Stream_23___mmap_RLAST;
  wire m_axi_rmem23___Mmap2Stream_23___mmap_RREADY;
  wire [1:0] m_axi_rmem23___Mmap2Stream_23___mmap_RRESP;
  wire m_axi_rmem23___Mmap2Stream_23___mmap_RVALID;
  wire [511:0] m_axi_rmem23___Mmap2Stream_23___mmap_WDATA;
  wire m_axi_rmem23___Mmap2Stream_23___mmap_WLAST;
  wire m_axi_rmem23___Mmap2Stream_23___mmap_WREADY;
  wire [63:0] m_axi_rmem23___Mmap2Stream_23___mmap_WSTRB;
  wire m_axi_rmem23___Mmap2Stream_23___mmap_WVALID;
  wire [63:0] m_axi_rmem23___Stream2Mmap_23___mmap_ARADDR;
  wire [1:0] m_axi_rmem23___Stream2Mmap_23___mmap_ARBURST;
  wire [3:0] m_axi_rmem23___Stream2Mmap_23___mmap_ARCACHE;
  wire [0:0] m_axi_rmem23___Stream2Mmap_23___mmap_ARID;
  wire [7:0] m_axi_rmem23___Stream2Mmap_23___mmap_ARLEN;
  wire m_axi_rmem23___Stream2Mmap_23___mmap_ARLOCK;
  wire [2:0] m_axi_rmem23___Stream2Mmap_23___mmap_ARPROT;
  wire [3:0] m_axi_rmem23___Stream2Mmap_23___mmap_ARQOS;
  wire m_axi_rmem23___Stream2Mmap_23___mmap_ARREADY;
  wire [2:0] m_axi_rmem23___Stream2Mmap_23___mmap_ARSIZE;
  wire m_axi_rmem23___Stream2Mmap_23___mmap_ARVALID;
  wire [63:0] m_axi_rmem23___Stream2Mmap_23___mmap_AWADDR;
  wire [1:0] m_axi_rmem23___Stream2Mmap_23___mmap_AWBURST;
  wire [3:0] m_axi_rmem23___Stream2Mmap_23___mmap_AWCACHE;
  wire [0:0] m_axi_rmem23___Stream2Mmap_23___mmap_AWID;
  wire [7:0] m_axi_rmem23___Stream2Mmap_23___mmap_AWLEN;
  wire m_axi_rmem23___Stream2Mmap_23___mmap_AWLOCK;
  wire [2:0] m_axi_rmem23___Stream2Mmap_23___mmap_AWPROT;
  wire [3:0] m_axi_rmem23___Stream2Mmap_23___mmap_AWQOS;
  wire m_axi_rmem23___Stream2Mmap_23___mmap_AWREADY;
  wire [2:0] m_axi_rmem23___Stream2Mmap_23___mmap_AWSIZE;
  wire m_axi_rmem23___Stream2Mmap_23___mmap_AWVALID;
  wire [0:0] m_axi_rmem23___Stream2Mmap_23___mmap_BID;
  wire m_axi_rmem23___Stream2Mmap_23___mmap_BREADY;
  wire [1:0] m_axi_rmem23___Stream2Mmap_23___mmap_BRESP;
  wire m_axi_rmem23___Stream2Mmap_23___mmap_BVALID;
  wire [511:0] m_axi_rmem23___Stream2Mmap_23___mmap_RDATA;
  wire [0:0] m_axi_rmem23___Stream2Mmap_23___mmap_RID;
  wire m_axi_rmem23___Stream2Mmap_23___mmap_RLAST;
  wire m_axi_rmem23___Stream2Mmap_23___mmap_RREADY;
  wire [1:0] m_axi_rmem23___Stream2Mmap_23___mmap_RRESP;
  wire m_axi_rmem23___Stream2Mmap_23___mmap_RVALID;
  wire [511:0] m_axi_rmem23___Stream2Mmap_23___mmap_WDATA;
  wire m_axi_rmem23___Stream2Mmap_23___mmap_WLAST;
  wire m_axi_rmem23___Stream2Mmap_23___mmap_WREADY;
  wire [63:0] m_axi_rmem23___Stream2Mmap_23___mmap_WSTRB;
  wire m_axi_rmem23___Stream2Mmap_23___mmap_WVALID;
  wire [63:0] m_axi_rmem24___Mmap2Stream_24___mmap_ARADDR;
  wire [1:0] m_axi_rmem24___Mmap2Stream_24___mmap_ARBURST;
  wire [3:0] m_axi_rmem24___Mmap2Stream_24___mmap_ARCACHE;
  wire [0:0] m_axi_rmem24___Mmap2Stream_24___mmap_ARID;
  wire [7:0] m_axi_rmem24___Mmap2Stream_24___mmap_ARLEN;
  wire m_axi_rmem24___Mmap2Stream_24___mmap_ARLOCK;
  wire [2:0] m_axi_rmem24___Mmap2Stream_24___mmap_ARPROT;
  wire [3:0] m_axi_rmem24___Mmap2Stream_24___mmap_ARQOS;
  wire m_axi_rmem24___Mmap2Stream_24___mmap_ARREADY;
  wire [2:0] m_axi_rmem24___Mmap2Stream_24___mmap_ARSIZE;
  wire m_axi_rmem24___Mmap2Stream_24___mmap_ARVALID;
  wire [63:0] m_axi_rmem24___Mmap2Stream_24___mmap_AWADDR;
  wire [1:0] m_axi_rmem24___Mmap2Stream_24___mmap_AWBURST;
  wire [3:0] m_axi_rmem24___Mmap2Stream_24___mmap_AWCACHE;
  wire [0:0] m_axi_rmem24___Mmap2Stream_24___mmap_AWID;
  wire [7:0] m_axi_rmem24___Mmap2Stream_24___mmap_AWLEN;
  wire m_axi_rmem24___Mmap2Stream_24___mmap_AWLOCK;
  wire [2:0] m_axi_rmem24___Mmap2Stream_24___mmap_AWPROT;
  wire [3:0] m_axi_rmem24___Mmap2Stream_24___mmap_AWQOS;
  wire m_axi_rmem24___Mmap2Stream_24___mmap_AWREADY;
  wire [2:0] m_axi_rmem24___Mmap2Stream_24___mmap_AWSIZE;
  wire m_axi_rmem24___Mmap2Stream_24___mmap_AWVALID;
  wire [0:0] m_axi_rmem24___Mmap2Stream_24___mmap_BID;
  wire m_axi_rmem24___Mmap2Stream_24___mmap_BREADY;
  wire [1:0] m_axi_rmem24___Mmap2Stream_24___mmap_BRESP;
  wire m_axi_rmem24___Mmap2Stream_24___mmap_BVALID;
  wire [511:0] m_axi_rmem24___Mmap2Stream_24___mmap_RDATA;
  wire [0:0] m_axi_rmem24___Mmap2Stream_24___mmap_RID;
  wire m_axi_rmem24___Mmap2Stream_24___mmap_RLAST;
  wire m_axi_rmem24___Mmap2Stream_24___mmap_RREADY;
  wire [1:0] m_axi_rmem24___Mmap2Stream_24___mmap_RRESP;
  wire m_axi_rmem24___Mmap2Stream_24___mmap_RVALID;
  wire [511:0] m_axi_rmem24___Mmap2Stream_24___mmap_WDATA;
  wire m_axi_rmem24___Mmap2Stream_24___mmap_WLAST;
  wire m_axi_rmem24___Mmap2Stream_24___mmap_WREADY;
  wire [63:0] m_axi_rmem24___Mmap2Stream_24___mmap_WSTRB;
  wire m_axi_rmem24___Mmap2Stream_24___mmap_WVALID;
  wire [63:0] m_axi_rmem24___Stream2Mmap_24___mmap_ARADDR;
  wire [1:0] m_axi_rmem24___Stream2Mmap_24___mmap_ARBURST;
  wire [3:0] m_axi_rmem24___Stream2Mmap_24___mmap_ARCACHE;
  wire [0:0] m_axi_rmem24___Stream2Mmap_24___mmap_ARID;
  wire [7:0] m_axi_rmem24___Stream2Mmap_24___mmap_ARLEN;
  wire m_axi_rmem24___Stream2Mmap_24___mmap_ARLOCK;
  wire [2:0] m_axi_rmem24___Stream2Mmap_24___mmap_ARPROT;
  wire [3:0] m_axi_rmem24___Stream2Mmap_24___mmap_ARQOS;
  wire m_axi_rmem24___Stream2Mmap_24___mmap_ARREADY;
  wire [2:0] m_axi_rmem24___Stream2Mmap_24___mmap_ARSIZE;
  wire m_axi_rmem24___Stream2Mmap_24___mmap_ARVALID;
  wire [63:0] m_axi_rmem24___Stream2Mmap_24___mmap_AWADDR;
  wire [1:0] m_axi_rmem24___Stream2Mmap_24___mmap_AWBURST;
  wire [3:0] m_axi_rmem24___Stream2Mmap_24___mmap_AWCACHE;
  wire [0:0] m_axi_rmem24___Stream2Mmap_24___mmap_AWID;
  wire [7:0] m_axi_rmem24___Stream2Mmap_24___mmap_AWLEN;
  wire m_axi_rmem24___Stream2Mmap_24___mmap_AWLOCK;
  wire [2:0] m_axi_rmem24___Stream2Mmap_24___mmap_AWPROT;
  wire [3:0] m_axi_rmem24___Stream2Mmap_24___mmap_AWQOS;
  wire m_axi_rmem24___Stream2Mmap_24___mmap_AWREADY;
  wire [2:0] m_axi_rmem24___Stream2Mmap_24___mmap_AWSIZE;
  wire m_axi_rmem24___Stream2Mmap_24___mmap_AWVALID;
  wire [0:0] m_axi_rmem24___Stream2Mmap_24___mmap_BID;
  wire m_axi_rmem24___Stream2Mmap_24___mmap_BREADY;
  wire [1:0] m_axi_rmem24___Stream2Mmap_24___mmap_BRESP;
  wire m_axi_rmem24___Stream2Mmap_24___mmap_BVALID;
  wire [511:0] m_axi_rmem24___Stream2Mmap_24___mmap_RDATA;
  wire [0:0] m_axi_rmem24___Stream2Mmap_24___mmap_RID;
  wire m_axi_rmem24___Stream2Mmap_24___mmap_RLAST;
  wire m_axi_rmem24___Stream2Mmap_24___mmap_RREADY;
  wire [1:0] m_axi_rmem24___Stream2Mmap_24___mmap_RRESP;
  wire m_axi_rmem24___Stream2Mmap_24___mmap_RVALID;
  wire [511:0] m_axi_rmem24___Stream2Mmap_24___mmap_WDATA;
  wire m_axi_rmem24___Stream2Mmap_24___mmap_WLAST;
  wire m_axi_rmem24___Stream2Mmap_24___mmap_WREADY;
  wire [63:0] m_axi_rmem24___Stream2Mmap_24___mmap_WSTRB;
  wire m_axi_rmem24___Stream2Mmap_24___mmap_WVALID;
  wire [63:0] m_axi_rmem25___Mmap2Stream_25___mmap_ARADDR;
  wire [1:0] m_axi_rmem25___Mmap2Stream_25___mmap_ARBURST;
  wire [3:0] m_axi_rmem25___Mmap2Stream_25___mmap_ARCACHE;
  wire [0:0] m_axi_rmem25___Mmap2Stream_25___mmap_ARID;
  wire [7:0] m_axi_rmem25___Mmap2Stream_25___mmap_ARLEN;
  wire m_axi_rmem25___Mmap2Stream_25___mmap_ARLOCK;
  wire [2:0] m_axi_rmem25___Mmap2Stream_25___mmap_ARPROT;
  wire [3:0] m_axi_rmem25___Mmap2Stream_25___mmap_ARQOS;
  wire m_axi_rmem25___Mmap2Stream_25___mmap_ARREADY;
  wire [2:0] m_axi_rmem25___Mmap2Stream_25___mmap_ARSIZE;
  wire m_axi_rmem25___Mmap2Stream_25___mmap_ARVALID;
  wire [63:0] m_axi_rmem25___Mmap2Stream_25___mmap_AWADDR;
  wire [1:0] m_axi_rmem25___Mmap2Stream_25___mmap_AWBURST;
  wire [3:0] m_axi_rmem25___Mmap2Stream_25___mmap_AWCACHE;
  wire [0:0] m_axi_rmem25___Mmap2Stream_25___mmap_AWID;
  wire [7:0] m_axi_rmem25___Mmap2Stream_25___mmap_AWLEN;
  wire m_axi_rmem25___Mmap2Stream_25___mmap_AWLOCK;
  wire [2:0] m_axi_rmem25___Mmap2Stream_25___mmap_AWPROT;
  wire [3:0] m_axi_rmem25___Mmap2Stream_25___mmap_AWQOS;
  wire m_axi_rmem25___Mmap2Stream_25___mmap_AWREADY;
  wire [2:0] m_axi_rmem25___Mmap2Stream_25___mmap_AWSIZE;
  wire m_axi_rmem25___Mmap2Stream_25___mmap_AWVALID;
  wire [0:0] m_axi_rmem25___Mmap2Stream_25___mmap_BID;
  wire m_axi_rmem25___Mmap2Stream_25___mmap_BREADY;
  wire [1:0] m_axi_rmem25___Mmap2Stream_25___mmap_BRESP;
  wire m_axi_rmem25___Mmap2Stream_25___mmap_BVALID;
  wire [511:0] m_axi_rmem25___Mmap2Stream_25___mmap_RDATA;
  wire [0:0] m_axi_rmem25___Mmap2Stream_25___mmap_RID;
  wire m_axi_rmem25___Mmap2Stream_25___mmap_RLAST;
  wire m_axi_rmem25___Mmap2Stream_25___mmap_RREADY;
  wire [1:0] m_axi_rmem25___Mmap2Stream_25___mmap_RRESP;
  wire m_axi_rmem25___Mmap2Stream_25___mmap_RVALID;
  wire [511:0] m_axi_rmem25___Mmap2Stream_25___mmap_WDATA;
  wire m_axi_rmem25___Mmap2Stream_25___mmap_WLAST;
  wire m_axi_rmem25___Mmap2Stream_25___mmap_WREADY;
  wire [63:0] m_axi_rmem25___Mmap2Stream_25___mmap_WSTRB;
  wire m_axi_rmem25___Mmap2Stream_25___mmap_WVALID;
  wire [63:0] m_axi_rmem25___Stream2Mmap_25___mmap_ARADDR;
  wire [1:0] m_axi_rmem25___Stream2Mmap_25___mmap_ARBURST;
  wire [3:0] m_axi_rmem25___Stream2Mmap_25___mmap_ARCACHE;
  wire [0:0] m_axi_rmem25___Stream2Mmap_25___mmap_ARID;
  wire [7:0] m_axi_rmem25___Stream2Mmap_25___mmap_ARLEN;
  wire m_axi_rmem25___Stream2Mmap_25___mmap_ARLOCK;
  wire [2:0] m_axi_rmem25___Stream2Mmap_25___mmap_ARPROT;
  wire [3:0] m_axi_rmem25___Stream2Mmap_25___mmap_ARQOS;
  wire m_axi_rmem25___Stream2Mmap_25___mmap_ARREADY;
  wire [2:0] m_axi_rmem25___Stream2Mmap_25___mmap_ARSIZE;
  wire m_axi_rmem25___Stream2Mmap_25___mmap_ARVALID;
  wire [63:0] m_axi_rmem25___Stream2Mmap_25___mmap_AWADDR;
  wire [1:0] m_axi_rmem25___Stream2Mmap_25___mmap_AWBURST;
  wire [3:0] m_axi_rmem25___Stream2Mmap_25___mmap_AWCACHE;
  wire [0:0] m_axi_rmem25___Stream2Mmap_25___mmap_AWID;
  wire [7:0] m_axi_rmem25___Stream2Mmap_25___mmap_AWLEN;
  wire m_axi_rmem25___Stream2Mmap_25___mmap_AWLOCK;
  wire [2:0] m_axi_rmem25___Stream2Mmap_25___mmap_AWPROT;
  wire [3:0] m_axi_rmem25___Stream2Mmap_25___mmap_AWQOS;
  wire m_axi_rmem25___Stream2Mmap_25___mmap_AWREADY;
  wire [2:0] m_axi_rmem25___Stream2Mmap_25___mmap_AWSIZE;
  wire m_axi_rmem25___Stream2Mmap_25___mmap_AWVALID;
  wire [0:0] m_axi_rmem25___Stream2Mmap_25___mmap_BID;
  wire m_axi_rmem25___Stream2Mmap_25___mmap_BREADY;
  wire [1:0] m_axi_rmem25___Stream2Mmap_25___mmap_BRESP;
  wire m_axi_rmem25___Stream2Mmap_25___mmap_BVALID;
  wire [511:0] m_axi_rmem25___Stream2Mmap_25___mmap_RDATA;
  wire [0:0] m_axi_rmem25___Stream2Mmap_25___mmap_RID;
  wire m_axi_rmem25___Stream2Mmap_25___mmap_RLAST;
  wire m_axi_rmem25___Stream2Mmap_25___mmap_RREADY;
  wire [1:0] m_axi_rmem25___Stream2Mmap_25___mmap_RRESP;
  wire m_axi_rmem25___Stream2Mmap_25___mmap_RVALID;
  wire [511:0] m_axi_rmem25___Stream2Mmap_25___mmap_WDATA;
  wire m_axi_rmem25___Stream2Mmap_25___mmap_WLAST;
  wire m_axi_rmem25___Stream2Mmap_25___mmap_WREADY;
  wire [63:0] m_axi_rmem25___Stream2Mmap_25___mmap_WSTRB;
  wire m_axi_rmem25___Stream2Mmap_25___mmap_WVALID;
  wire [63:0] m_axi_rmem26___Mmap2Stream_26___mmap_ARADDR;
  wire [1:0] m_axi_rmem26___Mmap2Stream_26___mmap_ARBURST;
  wire [3:0] m_axi_rmem26___Mmap2Stream_26___mmap_ARCACHE;
  wire [0:0] m_axi_rmem26___Mmap2Stream_26___mmap_ARID;
  wire [7:0] m_axi_rmem26___Mmap2Stream_26___mmap_ARLEN;
  wire m_axi_rmem26___Mmap2Stream_26___mmap_ARLOCK;
  wire [2:0] m_axi_rmem26___Mmap2Stream_26___mmap_ARPROT;
  wire [3:0] m_axi_rmem26___Mmap2Stream_26___mmap_ARQOS;
  wire m_axi_rmem26___Mmap2Stream_26___mmap_ARREADY;
  wire [2:0] m_axi_rmem26___Mmap2Stream_26___mmap_ARSIZE;
  wire m_axi_rmem26___Mmap2Stream_26___mmap_ARVALID;
  wire [63:0] m_axi_rmem26___Mmap2Stream_26___mmap_AWADDR;
  wire [1:0] m_axi_rmem26___Mmap2Stream_26___mmap_AWBURST;
  wire [3:0] m_axi_rmem26___Mmap2Stream_26___mmap_AWCACHE;
  wire [0:0] m_axi_rmem26___Mmap2Stream_26___mmap_AWID;
  wire [7:0] m_axi_rmem26___Mmap2Stream_26___mmap_AWLEN;
  wire m_axi_rmem26___Mmap2Stream_26___mmap_AWLOCK;
  wire [2:0] m_axi_rmem26___Mmap2Stream_26___mmap_AWPROT;
  wire [3:0] m_axi_rmem26___Mmap2Stream_26___mmap_AWQOS;
  wire m_axi_rmem26___Mmap2Stream_26___mmap_AWREADY;
  wire [2:0] m_axi_rmem26___Mmap2Stream_26___mmap_AWSIZE;
  wire m_axi_rmem26___Mmap2Stream_26___mmap_AWVALID;
  wire [0:0] m_axi_rmem26___Mmap2Stream_26___mmap_BID;
  wire m_axi_rmem26___Mmap2Stream_26___mmap_BREADY;
  wire [1:0] m_axi_rmem26___Mmap2Stream_26___mmap_BRESP;
  wire m_axi_rmem26___Mmap2Stream_26___mmap_BVALID;
  wire [511:0] m_axi_rmem26___Mmap2Stream_26___mmap_RDATA;
  wire [0:0] m_axi_rmem26___Mmap2Stream_26___mmap_RID;
  wire m_axi_rmem26___Mmap2Stream_26___mmap_RLAST;
  wire m_axi_rmem26___Mmap2Stream_26___mmap_RREADY;
  wire [1:0] m_axi_rmem26___Mmap2Stream_26___mmap_RRESP;
  wire m_axi_rmem26___Mmap2Stream_26___mmap_RVALID;
  wire [511:0] m_axi_rmem26___Mmap2Stream_26___mmap_WDATA;
  wire m_axi_rmem26___Mmap2Stream_26___mmap_WLAST;
  wire m_axi_rmem26___Mmap2Stream_26___mmap_WREADY;
  wire [63:0] m_axi_rmem26___Mmap2Stream_26___mmap_WSTRB;
  wire m_axi_rmem26___Mmap2Stream_26___mmap_WVALID;
  wire [63:0] m_axi_rmem26___Stream2Mmap_26___mmap_ARADDR;
  wire [1:0] m_axi_rmem26___Stream2Mmap_26___mmap_ARBURST;
  wire [3:0] m_axi_rmem26___Stream2Mmap_26___mmap_ARCACHE;
  wire [0:0] m_axi_rmem26___Stream2Mmap_26___mmap_ARID;
  wire [7:0] m_axi_rmem26___Stream2Mmap_26___mmap_ARLEN;
  wire m_axi_rmem26___Stream2Mmap_26___mmap_ARLOCK;
  wire [2:0] m_axi_rmem26___Stream2Mmap_26___mmap_ARPROT;
  wire [3:0] m_axi_rmem26___Stream2Mmap_26___mmap_ARQOS;
  wire m_axi_rmem26___Stream2Mmap_26___mmap_ARREADY;
  wire [2:0] m_axi_rmem26___Stream2Mmap_26___mmap_ARSIZE;
  wire m_axi_rmem26___Stream2Mmap_26___mmap_ARVALID;
  wire [63:0] m_axi_rmem26___Stream2Mmap_26___mmap_AWADDR;
  wire [1:0] m_axi_rmem26___Stream2Mmap_26___mmap_AWBURST;
  wire [3:0] m_axi_rmem26___Stream2Mmap_26___mmap_AWCACHE;
  wire [0:0] m_axi_rmem26___Stream2Mmap_26___mmap_AWID;
  wire [7:0] m_axi_rmem26___Stream2Mmap_26___mmap_AWLEN;
  wire m_axi_rmem26___Stream2Mmap_26___mmap_AWLOCK;
  wire [2:0] m_axi_rmem26___Stream2Mmap_26___mmap_AWPROT;
  wire [3:0] m_axi_rmem26___Stream2Mmap_26___mmap_AWQOS;
  wire m_axi_rmem26___Stream2Mmap_26___mmap_AWREADY;
  wire [2:0] m_axi_rmem26___Stream2Mmap_26___mmap_AWSIZE;
  wire m_axi_rmem26___Stream2Mmap_26___mmap_AWVALID;
  wire [0:0] m_axi_rmem26___Stream2Mmap_26___mmap_BID;
  wire m_axi_rmem26___Stream2Mmap_26___mmap_BREADY;
  wire [1:0] m_axi_rmem26___Stream2Mmap_26___mmap_BRESP;
  wire m_axi_rmem26___Stream2Mmap_26___mmap_BVALID;
  wire [511:0] m_axi_rmem26___Stream2Mmap_26___mmap_RDATA;
  wire [0:0] m_axi_rmem26___Stream2Mmap_26___mmap_RID;
  wire m_axi_rmem26___Stream2Mmap_26___mmap_RLAST;
  wire m_axi_rmem26___Stream2Mmap_26___mmap_RREADY;
  wire [1:0] m_axi_rmem26___Stream2Mmap_26___mmap_RRESP;
  wire m_axi_rmem26___Stream2Mmap_26___mmap_RVALID;
  wire [511:0] m_axi_rmem26___Stream2Mmap_26___mmap_WDATA;
  wire m_axi_rmem26___Stream2Mmap_26___mmap_WLAST;
  wire m_axi_rmem26___Stream2Mmap_26___mmap_WREADY;
  wire [63:0] m_axi_rmem26___Stream2Mmap_26___mmap_WSTRB;
  wire m_axi_rmem26___Stream2Mmap_26___mmap_WVALID;
  wire [63:0] m_axi_rmem27___Mmap2Stream_27___mmap_ARADDR;
  wire [1:0] m_axi_rmem27___Mmap2Stream_27___mmap_ARBURST;
  wire [3:0] m_axi_rmem27___Mmap2Stream_27___mmap_ARCACHE;
  wire [0:0] m_axi_rmem27___Mmap2Stream_27___mmap_ARID;
  wire [7:0] m_axi_rmem27___Mmap2Stream_27___mmap_ARLEN;
  wire m_axi_rmem27___Mmap2Stream_27___mmap_ARLOCK;
  wire [2:0] m_axi_rmem27___Mmap2Stream_27___mmap_ARPROT;
  wire [3:0] m_axi_rmem27___Mmap2Stream_27___mmap_ARQOS;
  wire m_axi_rmem27___Mmap2Stream_27___mmap_ARREADY;
  wire [2:0] m_axi_rmem27___Mmap2Stream_27___mmap_ARSIZE;
  wire m_axi_rmem27___Mmap2Stream_27___mmap_ARVALID;
  wire [63:0] m_axi_rmem27___Mmap2Stream_27___mmap_AWADDR;
  wire [1:0] m_axi_rmem27___Mmap2Stream_27___mmap_AWBURST;
  wire [3:0] m_axi_rmem27___Mmap2Stream_27___mmap_AWCACHE;
  wire [0:0] m_axi_rmem27___Mmap2Stream_27___mmap_AWID;
  wire [7:0] m_axi_rmem27___Mmap2Stream_27___mmap_AWLEN;
  wire m_axi_rmem27___Mmap2Stream_27___mmap_AWLOCK;
  wire [2:0] m_axi_rmem27___Mmap2Stream_27___mmap_AWPROT;
  wire [3:0] m_axi_rmem27___Mmap2Stream_27___mmap_AWQOS;
  wire m_axi_rmem27___Mmap2Stream_27___mmap_AWREADY;
  wire [2:0] m_axi_rmem27___Mmap2Stream_27___mmap_AWSIZE;
  wire m_axi_rmem27___Mmap2Stream_27___mmap_AWVALID;
  wire [0:0] m_axi_rmem27___Mmap2Stream_27___mmap_BID;
  wire m_axi_rmem27___Mmap2Stream_27___mmap_BREADY;
  wire [1:0] m_axi_rmem27___Mmap2Stream_27___mmap_BRESP;
  wire m_axi_rmem27___Mmap2Stream_27___mmap_BVALID;
  wire [511:0] m_axi_rmem27___Mmap2Stream_27___mmap_RDATA;
  wire [0:0] m_axi_rmem27___Mmap2Stream_27___mmap_RID;
  wire m_axi_rmem27___Mmap2Stream_27___mmap_RLAST;
  wire m_axi_rmem27___Mmap2Stream_27___mmap_RREADY;
  wire [1:0] m_axi_rmem27___Mmap2Stream_27___mmap_RRESP;
  wire m_axi_rmem27___Mmap2Stream_27___mmap_RVALID;
  wire [511:0] m_axi_rmem27___Mmap2Stream_27___mmap_WDATA;
  wire m_axi_rmem27___Mmap2Stream_27___mmap_WLAST;
  wire m_axi_rmem27___Mmap2Stream_27___mmap_WREADY;
  wire [63:0] m_axi_rmem27___Mmap2Stream_27___mmap_WSTRB;
  wire m_axi_rmem27___Mmap2Stream_27___mmap_WVALID;
  wire [63:0] m_axi_rmem27___Stream2Mmap_27___mmap_ARADDR;
  wire [1:0] m_axi_rmem27___Stream2Mmap_27___mmap_ARBURST;
  wire [3:0] m_axi_rmem27___Stream2Mmap_27___mmap_ARCACHE;
  wire [0:0] m_axi_rmem27___Stream2Mmap_27___mmap_ARID;
  wire [7:0] m_axi_rmem27___Stream2Mmap_27___mmap_ARLEN;
  wire m_axi_rmem27___Stream2Mmap_27___mmap_ARLOCK;
  wire [2:0] m_axi_rmem27___Stream2Mmap_27___mmap_ARPROT;
  wire [3:0] m_axi_rmem27___Stream2Mmap_27___mmap_ARQOS;
  wire m_axi_rmem27___Stream2Mmap_27___mmap_ARREADY;
  wire [2:0] m_axi_rmem27___Stream2Mmap_27___mmap_ARSIZE;
  wire m_axi_rmem27___Stream2Mmap_27___mmap_ARVALID;
  wire [63:0] m_axi_rmem27___Stream2Mmap_27___mmap_AWADDR;
  wire [1:0] m_axi_rmem27___Stream2Mmap_27___mmap_AWBURST;
  wire [3:0] m_axi_rmem27___Stream2Mmap_27___mmap_AWCACHE;
  wire [0:0] m_axi_rmem27___Stream2Mmap_27___mmap_AWID;
  wire [7:0] m_axi_rmem27___Stream2Mmap_27___mmap_AWLEN;
  wire m_axi_rmem27___Stream2Mmap_27___mmap_AWLOCK;
  wire [2:0] m_axi_rmem27___Stream2Mmap_27___mmap_AWPROT;
  wire [3:0] m_axi_rmem27___Stream2Mmap_27___mmap_AWQOS;
  wire m_axi_rmem27___Stream2Mmap_27___mmap_AWREADY;
  wire [2:0] m_axi_rmem27___Stream2Mmap_27___mmap_AWSIZE;
  wire m_axi_rmem27___Stream2Mmap_27___mmap_AWVALID;
  wire [0:0] m_axi_rmem27___Stream2Mmap_27___mmap_BID;
  wire m_axi_rmem27___Stream2Mmap_27___mmap_BREADY;
  wire [1:0] m_axi_rmem27___Stream2Mmap_27___mmap_BRESP;
  wire m_axi_rmem27___Stream2Mmap_27___mmap_BVALID;
  wire [511:0] m_axi_rmem27___Stream2Mmap_27___mmap_RDATA;
  wire [0:0] m_axi_rmem27___Stream2Mmap_27___mmap_RID;
  wire m_axi_rmem27___Stream2Mmap_27___mmap_RLAST;
  wire m_axi_rmem27___Stream2Mmap_27___mmap_RREADY;
  wire [1:0] m_axi_rmem27___Stream2Mmap_27___mmap_RRESP;
  wire m_axi_rmem27___Stream2Mmap_27___mmap_RVALID;
  wire [511:0] m_axi_rmem27___Stream2Mmap_27___mmap_WDATA;
  wire m_axi_rmem27___Stream2Mmap_27___mmap_WLAST;
  wire m_axi_rmem27___Stream2Mmap_27___mmap_WREADY;
  wire [63:0] m_axi_rmem27___Stream2Mmap_27___mmap_WSTRB;
  wire m_axi_rmem27___Stream2Mmap_27___mmap_WVALID;
  wire [63:0] Mmap2Stream_0___n__q0;
  wire [63:0] Mmap2Stream_0___rmem0__q0;
  wire Mmap2Stream_0__ap_start;
  wire Mmap2Stream_0__ap_ready;
  wire Mmap2Stream_0__ap_done;
  wire Mmap2Stream_0__ap_idle;
  wire [63:0] Mmap2Stream_1___n__q0;
  wire [63:0] Mmap2Stream_1___rmem1__q0;
  wire Mmap2Stream_1__ap_start;
  wire Mmap2Stream_1__ap_ready;
  wire Mmap2Stream_1__ap_done;
  wire Mmap2Stream_1__ap_idle;
  wire [63:0] Mmap2Stream_2___n__q0;
  wire [63:0] Mmap2Stream_2___rmem2__q0;
  wire Mmap2Stream_2__ap_start;
  wire Mmap2Stream_2__ap_ready;
  wire Mmap2Stream_2__ap_done;
  wire Mmap2Stream_2__ap_idle;
  wire [63:0] Mmap2Stream_3___n__q0;
  wire [63:0] Mmap2Stream_3___rmem3__q0;
  wire Mmap2Stream_3__ap_start;
  wire Mmap2Stream_3__ap_ready;
  wire Mmap2Stream_3__ap_done;
  wire Mmap2Stream_3__ap_idle;
  wire [63:0] Mmap2Stream_4___n__q0;
  wire [63:0] Mmap2Stream_4___rmem4__q0;
  wire Mmap2Stream_4__ap_start;
  wire Mmap2Stream_4__ap_ready;
  wire Mmap2Stream_4__ap_done;
  wire Mmap2Stream_4__ap_idle;
  wire [63:0] Mmap2Stream_5___n__q0;
  wire [63:0] Mmap2Stream_5___rmem5__q0;
  wire Mmap2Stream_5__ap_start;
  wire Mmap2Stream_5__ap_ready;
  wire Mmap2Stream_5__ap_done;
  wire Mmap2Stream_5__ap_idle;
  wire [63:0] Mmap2Stream_6___n__q0;
  wire [63:0] Mmap2Stream_6___rmem6__q0;
  wire Mmap2Stream_6__ap_start;
  wire Mmap2Stream_6__ap_ready;
  wire Mmap2Stream_6__ap_done;
  wire Mmap2Stream_6__ap_idle;
  wire [63:0] Mmap2Stream_7___n__q0;
  wire [63:0] Mmap2Stream_7___rmem7__q0;
  wire Mmap2Stream_7__ap_start;
  wire Mmap2Stream_7__ap_ready;
  wire Mmap2Stream_7__ap_done;
  wire Mmap2Stream_7__ap_idle;
  wire [63:0] Mmap2Stream_8___n__q0;
  wire [63:0] Mmap2Stream_8___rmem8__q0;
  wire Mmap2Stream_8__ap_start;
  wire Mmap2Stream_8__ap_ready;
  wire Mmap2Stream_8__ap_done;
  wire Mmap2Stream_8__ap_idle;
  wire [63:0] Mmap2Stream_9___n__q0;
  wire [63:0] Mmap2Stream_9___rmem9__q0;
  wire Mmap2Stream_9__ap_start;
  wire Mmap2Stream_9__ap_ready;
  wire Mmap2Stream_9__ap_done;
  wire Mmap2Stream_9__ap_idle;
  wire [63:0] Mmap2Stream_10___n__q0;
  wire [63:0] Mmap2Stream_10___rmem10__q0;
  wire Mmap2Stream_10__ap_start;
  wire Mmap2Stream_10__ap_ready;
  wire Mmap2Stream_10__ap_done;
  wire Mmap2Stream_10__ap_idle;
  wire [63:0] Mmap2Stream_11___n__q0;
  wire [63:0] Mmap2Stream_11___rmem11__q0;
  wire Mmap2Stream_11__ap_start;
  wire Mmap2Stream_11__ap_ready;
  wire Mmap2Stream_11__ap_done;
  wire Mmap2Stream_11__ap_idle;
  wire [63:0] Mmap2Stream_12___n__q0;
  wire [63:0] Mmap2Stream_12___rmem12__q0;
  wire Mmap2Stream_12__ap_start;
  wire Mmap2Stream_12__ap_ready;
  wire Mmap2Stream_12__ap_done;
  wire Mmap2Stream_12__ap_idle;
  wire [63:0] Mmap2Stream_13___n__q0;
  wire [63:0] Mmap2Stream_13___rmem13__q0;
  wire Mmap2Stream_13__ap_start;
  wire Mmap2Stream_13__ap_ready;
  wire Mmap2Stream_13__ap_done;
  wire Mmap2Stream_13__ap_idle;
  wire [63:0] Mmap2Stream_14___n__q0;
  wire [63:0] Mmap2Stream_14___rmem14__q0;
  wire Mmap2Stream_14__ap_start;
  wire Mmap2Stream_14__ap_ready;
  wire Mmap2Stream_14__ap_done;
  wire Mmap2Stream_14__ap_idle;
  wire [63:0] Mmap2Stream_15___n__q0;
  wire [63:0] Mmap2Stream_15___rmem15__q0;
  wire Mmap2Stream_15__ap_start;
  wire Mmap2Stream_15__ap_ready;
  wire Mmap2Stream_15__ap_done;
  wire Mmap2Stream_15__ap_idle;
  wire [63:0] Mmap2Stream_16___n__q0;
  wire [63:0] Mmap2Stream_16___rmem16__q0;
  wire Mmap2Stream_16__ap_start;
  wire Mmap2Stream_16__ap_ready;
  wire Mmap2Stream_16__ap_done;
  wire Mmap2Stream_16__ap_idle;
  wire [63:0] Mmap2Stream_17___n__q0;
  wire [63:0] Mmap2Stream_17___rmem17__q0;
  wire Mmap2Stream_17__ap_start;
  wire Mmap2Stream_17__ap_ready;
  wire Mmap2Stream_17__ap_done;
  wire Mmap2Stream_17__ap_idle;
  wire [63:0] Mmap2Stream_18___n__q0;
  wire [63:0] Mmap2Stream_18___rmem18__q0;
  wire Mmap2Stream_18__ap_start;
  wire Mmap2Stream_18__ap_ready;
  wire Mmap2Stream_18__ap_done;
  wire Mmap2Stream_18__ap_idle;
  wire [63:0] Mmap2Stream_19___n__q0;
  wire [63:0] Mmap2Stream_19___rmem19__q0;
  wire Mmap2Stream_19__ap_start;
  wire Mmap2Stream_19__ap_ready;
  wire Mmap2Stream_19__ap_done;
  wire Mmap2Stream_19__ap_idle;
  wire [63:0] Mmap2Stream_20___n__q0;
  wire [63:0] Mmap2Stream_20___rmem20__q0;
  wire Mmap2Stream_20__ap_start;
  wire Mmap2Stream_20__ap_ready;
  wire Mmap2Stream_20__ap_done;
  wire Mmap2Stream_20__ap_idle;
  wire [63:0] Mmap2Stream_21___n__q0;
  wire [63:0] Mmap2Stream_21___rmem21__q0;
  wire Mmap2Stream_21__ap_start;
  wire Mmap2Stream_21__ap_ready;
  wire Mmap2Stream_21__ap_done;
  wire Mmap2Stream_21__ap_idle;
  wire [63:0] Mmap2Stream_22___n__q0;
  wire [63:0] Mmap2Stream_22___rmem22__q0;
  wire Mmap2Stream_22__ap_start;
  wire Mmap2Stream_22__ap_ready;
  wire Mmap2Stream_22__ap_done;
  wire Mmap2Stream_22__ap_idle;
  wire [63:0] Mmap2Stream_23___n__q0;
  wire [63:0] Mmap2Stream_23___rmem23__q0;
  wire Mmap2Stream_23__ap_start;
  wire Mmap2Stream_23__ap_ready;
  wire Mmap2Stream_23__ap_done;
  wire Mmap2Stream_23__ap_idle;
  wire [63:0] Mmap2Stream_24___n__q0;
  wire [63:0] Mmap2Stream_24___rmem24__q0;
  wire Mmap2Stream_24__ap_start;
  wire Mmap2Stream_24__ap_ready;
  wire Mmap2Stream_24__ap_done;
  wire Mmap2Stream_24__ap_idle;
  wire [63:0] Mmap2Stream_25___n__q0;
  wire [63:0] Mmap2Stream_25___rmem25__q0;
  wire Mmap2Stream_25__ap_start;
  wire Mmap2Stream_25__ap_ready;
  wire Mmap2Stream_25__ap_done;
  wire Mmap2Stream_25__ap_idle;
  wire [63:0] Mmap2Stream_26___n__q0;
  wire [63:0] Mmap2Stream_26___rmem26__q0;
  wire Mmap2Stream_26__ap_start;
  wire Mmap2Stream_26__ap_ready;
  wire Mmap2Stream_26__ap_done;
  wire Mmap2Stream_26__ap_idle;
  wire [63:0] Mmap2Stream_27___n__q0;
  wire [63:0] Mmap2Stream_27___rmem27__q0;
  wire Mmap2Stream_27__ap_start;
  wire Mmap2Stream_27__ap_ready;
  wire Mmap2Stream_27__ap_done;
  wire Mmap2Stream_27__ap_idle;
  wire [63:0] Stream2Mmap_0___n__q0;
  wire [63:0] Stream2Mmap_0___rmem0__q0;
  wire Stream2Mmap_0__ap_start;
  wire Stream2Mmap_0__ap_ready;
  wire Stream2Mmap_0__ap_done;
  wire Stream2Mmap_0__ap_idle;
  wire [63:0] Stream2Mmap_1___n__q0;
  wire [63:0] Stream2Mmap_1___rmem1__q0;
  wire Stream2Mmap_1__ap_start;
  wire Stream2Mmap_1__ap_ready;
  wire Stream2Mmap_1__ap_done;
  wire Stream2Mmap_1__ap_idle;
  wire [63:0] Stream2Mmap_2___n__q0;
  wire [63:0] Stream2Mmap_2___rmem2__q0;
  wire Stream2Mmap_2__ap_start;
  wire Stream2Mmap_2__ap_ready;
  wire Stream2Mmap_2__ap_done;
  wire Stream2Mmap_2__ap_idle;
  wire [63:0] Stream2Mmap_3___n__q0;
  wire [63:0] Stream2Mmap_3___rmem3__q0;
  wire Stream2Mmap_3__ap_start;
  wire Stream2Mmap_3__ap_ready;
  wire Stream2Mmap_3__ap_done;
  wire Stream2Mmap_3__ap_idle;
  wire [63:0] Stream2Mmap_4___n__q0;
  wire [63:0] Stream2Mmap_4___rmem4__q0;
  wire Stream2Mmap_4__ap_start;
  wire Stream2Mmap_4__ap_ready;
  wire Stream2Mmap_4__ap_done;
  wire Stream2Mmap_4__ap_idle;
  wire [63:0] Stream2Mmap_5___n__q0;
  wire [63:0] Stream2Mmap_5___rmem5__q0;
  wire Stream2Mmap_5__ap_start;
  wire Stream2Mmap_5__ap_ready;
  wire Stream2Mmap_5__ap_done;
  wire Stream2Mmap_5__ap_idle;
  wire [63:0] Stream2Mmap_6___n__q0;
  wire [63:0] Stream2Mmap_6___rmem6__q0;
  wire Stream2Mmap_6__ap_start;
  wire Stream2Mmap_6__ap_ready;
  wire Stream2Mmap_6__ap_done;
  wire Stream2Mmap_6__ap_idle;
  wire [63:0] Stream2Mmap_7___n__q0;
  wire [63:0] Stream2Mmap_7___rmem7__q0;
  wire Stream2Mmap_7__ap_start;
  wire Stream2Mmap_7__ap_ready;
  wire Stream2Mmap_7__ap_done;
  wire Stream2Mmap_7__ap_idle;
  wire [63:0] Stream2Mmap_8___n__q0;
  wire [63:0] Stream2Mmap_8___rmem8__q0;
  wire Stream2Mmap_8__ap_start;
  wire Stream2Mmap_8__ap_ready;
  wire Stream2Mmap_8__ap_done;
  wire Stream2Mmap_8__ap_idle;
  wire [63:0] Stream2Mmap_9___n__q0;
  wire [63:0] Stream2Mmap_9___rmem9__q0;
  wire Stream2Mmap_9__ap_start;
  wire Stream2Mmap_9__ap_ready;
  wire Stream2Mmap_9__ap_done;
  wire Stream2Mmap_9__ap_idle;
  wire [63:0] Stream2Mmap_10___n__q0;
  wire [63:0] Stream2Mmap_10___rmem10__q0;
  wire Stream2Mmap_10__ap_start;
  wire Stream2Mmap_10__ap_ready;
  wire Stream2Mmap_10__ap_done;
  wire Stream2Mmap_10__ap_idle;
  wire [63:0] Stream2Mmap_11___n__q0;
  wire [63:0] Stream2Mmap_11___rmem11__q0;
  wire Stream2Mmap_11__ap_start;
  wire Stream2Mmap_11__ap_ready;
  wire Stream2Mmap_11__ap_done;
  wire Stream2Mmap_11__ap_idle;
  wire [63:0] Stream2Mmap_12___n__q0;
  wire [63:0] Stream2Mmap_12___rmem12__q0;
  wire Stream2Mmap_12__ap_start;
  wire Stream2Mmap_12__ap_ready;
  wire Stream2Mmap_12__ap_done;
  wire Stream2Mmap_12__ap_idle;
  wire [63:0] Stream2Mmap_13___n__q0;
  wire [63:0] Stream2Mmap_13___rmem13__q0;
  wire Stream2Mmap_13__ap_start;
  wire Stream2Mmap_13__ap_ready;
  wire Stream2Mmap_13__ap_done;
  wire Stream2Mmap_13__ap_idle;
  wire [63:0] Stream2Mmap_14___n__q0;
  wire [63:0] Stream2Mmap_14___rmem14__q0;
  wire Stream2Mmap_14__ap_start;
  wire Stream2Mmap_14__ap_ready;
  wire Stream2Mmap_14__ap_done;
  wire Stream2Mmap_14__ap_idle;
  wire [63:0] Stream2Mmap_15___n__q0;
  wire [63:0] Stream2Mmap_15___rmem15__q0;
  wire Stream2Mmap_15__ap_start;
  wire Stream2Mmap_15__ap_ready;
  wire Stream2Mmap_15__ap_done;
  wire Stream2Mmap_15__ap_idle;
  wire [63:0] Stream2Mmap_16___n__q0;
  wire [63:0] Stream2Mmap_16___rmem16__q0;
  wire Stream2Mmap_16__ap_start;
  wire Stream2Mmap_16__ap_ready;
  wire Stream2Mmap_16__ap_done;
  wire Stream2Mmap_16__ap_idle;
  wire [63:0] Stream2Mmap_17___n__q0;
  wire [63:0] Stream2Mmap_17___rmem17__q0;
  wire Stream2Mmap_17__ap_start;
  wire Stream2Mmap_17__ap_ready;
  wire Stream2Mmap_17__ap_done;
  wire Stream2Mmap_17__ap_idle;
  wire [63:0] Stream2Mmap_18___n__q0;
  wire [63:0] Stream2Mmap_18___rmem18__q0;
  wire Stream2Mmap_18__ap_start;
  wire Stream2Mmap_18__ap_ready;
  wire Stream2Mmap_18__ap_done;
  wire Stream2Mmap_18__ap_idle;
  wire [63:0] Stream2Mmap_19___n__q0;
  wire [63:0] Stream2Mmap_19___rmem19__q0;
  wire Stream2Mmap_19__ap_start;
  wire Stream2Mmap_19__ap_ready;
  wire Stream2Mmap_19__ap_done;
  wire Stream2Mmap_19__ap_idle;
  wire [63:0] Stream2Mmap_20___n__q0;
  wire [63:0] Stream2Mmap_20___rmem20__q0;
  wire Stream2Mmap_20__ap_start;
  wire Stream2Mmap_20__ap_ready;
  wire Stream2Mmap_20__ap_done;
  wire Stream2Mmap_20__ap_idle;
  wire [63:0] Stream2Mmap_21___n__q0;
  wire [63:0] Stream2Mmap_21___rmem21__q0;
  wire Stream2Mmap_21__ap_start;
  wire Stream2Mmap_21__ap_ready;
  wire Stream2Mmap_21__ap_done;
  wire Stream2Mmap_21__ap_idle;
  wire [63:0] Stream2Mmap_22___n__q0;
  wire [63:0] Stream2Mmap_22___rmem22__q0;
  wire Stream2Mmap_22__ap_start;
  wire Stream2Mmap_22__ap_ready;
  wire Stream2Mmap_22__ap_done;
  wire Stream2Mmap_22__ap_idle;
  wire [63:0] Stream2Mmap_23___n__q0;
  wire [63:0] Stream2Mmap_23___rmem23__q0;
  wire Stream2Mmap_23__ap_start;
  wire Stream2Mmap_23__ap_ready;
  wire Stream2Mmap_23__ap_done;
  wire Stream2Mmap_23__ap_idle;
  wire [63:0] Stream2Mmap_24___n__q0;
  wire [63:0] Stream2Mmap_24___rmem24__q0;
  wire Stream2Mmap_24__ap_start;
  wire Stream2Mmap_24__ap_ready;
  wire Stream2Mmap_24__ap_done;
  wire Stream2Mmap_24__ap_idle;
  wire [63:0] Stream2Mmap_25___n__q0;
  wire [63:0] Stream2Mmap_25___rmem25__q0;
  wire Stream2Mmap_25__ap_start;
  wire Stream2Mmap_25__ap_ready;
  wire Stream2Mmap_25__ap_done;
  wire Stream2Mmap_25__ap_idle;
  wire [63:0] Stream2Mmap_26___n__q0;
  wire [63:0] Stream2Mmap_26___rmem26__q0;
  wire Stream2Mmap_26__ap_start;
  wire Stream2Mmap_26__ap_ready;
  wire Stream2Mmap_26__ap_done;
  wire Stream2Mmap_26__ap_idle;
  wire [63:0] Stream2Mmap_27___n__q0;
  wire [63:0] Stream2Mmap_27___rmem27__q0;
  wire Stream2Mmap_27__ap_start;
  wire Stream2Mmap_27__ap_ready;
  wire Stream2Mmap_27__ap_done;
  wire Stream2Mmap_27__ap_idle;
  wire [63:0] yshift_0___n__q0;
  wire yshift_0__ap_start;
  wire yshift_0__ap_ready;
  wire yshift_0__ap_done;
  wire yshift_0__ap_idle;
  wire [63:0] yshift_1___n__q0;
  wire yshift_1__ap_start;
  wire yshift_1__ap_ready;
  wire yshift_1__ap_done;
  wire yshift_1__ap_idle;
  wire [63:0] yshift_2___n__q0;
  wire yshift_2__ap_start;
  wire yshift_2__ap_ready;
  wire yshift_2__ap_done;
  wire yshift_2__ap_idle;
  wire [63:0] yshift_3___n__q0;
  wire yshift_3__ap_start;
  wire yshift_3__ap_ready;
  wire yshift_3__ap_done;
  wire yshift_3__ap_idle;
  wire [63:0] yshift_4___n__q0;
  wire yshift_4__ap_start;
  wire yshift_4__ap_ready;
  wire yshift_4__ap_done;
  wire yshift_4__ap_idle;
  wire [63:0] yshift_5___n__q0;
  wire yshift_5__ap_start;
  wire yshift_5__ap_ready;
  wire yshift_5__ap_done;
  wire yshift_5__ap_idle;
  wire [63:0] yshift_6___n__q0;
  wire yshift_6__ap_start;
  wire yshift_6__ap_ready;
  wire yshift_6__ap_done;
  wire yshift_6__ap_idle;
  wire [63:0] yshift_7___n__q0;
  wire yshift_7__ap_start;
  wire yshift_7__ap_ready;
  wire yshift_7__ap_done;
  wire yshift_7__ap_idle;
  wire [63:0] yshift_8___n__q0;
  wire yshift_8__ap_start;
  wire yshift_8__ap_ready;
  wire yshift_8__ap_done;
  wire yshift_8__ap_idle;
  wire [63:0] yshift_9___n__q0;
  wire yshift_9__ap_start;
  wire yshift_9__ap_ready;
  wire yshift_9__ap_done;
  wire yshift_9__ap_idle;
  wire [63:0] yshift_10___n__q0;
  wire yshift_10__ap_start;
  wire yshift_10__ap_ready;
  wire yshift_10__ap_done;
  wire yshift_10__ap_idle;
  wire [63:0] yshift_11___n__q0;
  wire yshift_11__ap_start;
  wire yshift_11__ap_ready;
  wire yshift_11__ap_done;
  wire yshift_11__ap_idle;
  wire [63:0] yshift_12___n__q0;
  wire yshift_12__ap_start;
  wire yshift_12__ap_ready;
  wire yshift_12__ap_done;
  wire yshift_12__ap_idle;
  wire [63:0] yshift_13___n__q0;
  wire yshift_13__ap_start;
  wire yshift_13__ap_ready;
  wire yshift_13__ap_done;
  wire yshift_13__ap_idle;
  wire [63:0] yshift_14___n__q0;
  wire yshift_14__ap_start;
  wire yshift_14__ap_ready;
  wire yshift_14__ap_done;
  wire yshift_14__ap_idle;
  wire [63:0] yshift_15___n__q0;
  wire yshift_15__ap_start;
  wire yshift_15__ap_ready;
  wire yshift_15__ap_done;
  wire yshift_15__ap_idle;
  wire [63:0] yshift_16___n__q0;
  wire yshift_16__ap_start;
  wire yshift_16__ap_ready;
  wire yshift_16__ap_done;
  wire yshift_16__ap_idle;
  wire [63:0] yshift_17___n__q0;
  wire yshift_17__ap_start;
  wire yshift_17__ap_ready;
  wire yshift_17__ap_done;
  wire yshift_17__ap_idle;
  wire [63:0] yshift_18___n__q0;
  wire yshift_18__ap_start;
  wire yshift_18__ap_ready;
  wire yshift_18__ap_done;
  wire yshift_18__ap_idle;
  wire [63:0] yshift_19___n__q0;
  wire yshift_19__ap_start;
  wire yshift_19__ap_ready;
  wire yshift_19__ap_done;
  wire yshift_19__ap_idle;
  wire [63:0] yshift_20___n__q0;
  wire yshift_20__ap_start;
  wire yshift_20__ap_ready;
  wire yshift_20__ap_done;
  wire yshift_20__ap_idle;
  wire [63:0] yshift_21___n__q0;
  wire yshift_21__ap_start;
  wire yshift_21__ap_ready;
  wire yshift_21__ap_done;
  wire yshift_21__ap_idle;
  wire [63:0] yshift_22___n__q0;
  wire yshift_22__ap_start;
  wire yshift_22__ap_ready;
  wire yshift_22__ap_done;
  wire yshift_22__ap_idle;
  wire [63:0] yshift_23___n__q0;
  wire yshift_23__ap_start;
  wire yshift_23__ap_ready;
  wire yshift_23__ap_done;
  wire yshift_23__ap_idle;
  wire [63:0] yshift_24___n__q0;
  wire yshift_24__ap_start;
  wire yshift_24__ap_ready;
  wire yshift_24__ap_done;
  wire yshift_24__ap_idle;
  wire [63:0] yshift_25___n__q0;
  wire yshift_25__ap_start;
  wire yshift_25__ap_ready;
  wire yshift_25__ap_done;
  wire yshift_25__ap_idle;
  wire [63:0] yshift_26___n__q0;
  wire yshift_26__ap_start;
  wire yshift_26__ap_ready;
  wire yshift_26__ap_done;
  wire yshift_26__ap_idle;
  wire [63:0] yshift_27___n__q0;
  wire yshift_27__ap_start;
  wire yshift_27__ap_ready;
  wire yshift_27__ap_done;
  wire yshift_27__ap_idle;
  wire ap_rst_n_inv;
  wire ap_done;
  wire ap_idle;
  wire ap_ready;

  vadd_bw_control_s_axi
  #(
    .C_S_AXI_ADDR_WIDTH(C_S_AXI_CONTROL_ADDR_WIDTH),
    .C_S_AXI_DATA_WIDTH(C_S_AXI_CONTROL_DATA_WIDTH)
  )
  control_s_axi_U
  (
    .AWVALID(s_axi_control_AWVALID),
    .AWREADY(s_axi_control_AWREADY),
    .AWADDR(s_axi_control_AWADDR),
    .WVALID(s_axi_control_WVALID),
    .WREADY(s_axi_control_WREADY),
    .WDATA(s_axi_control_WDATA),
    .WSTRB(s_axi_control_WSTRB),
    .ARVALID(s_axi_control_ARVALID),
    .ARREADY(s_axi_control_ARREADY),
    .ARADDR(s_axi_control_ARADDR),
    .RVALID(s_axi_control_RVALID),
    .RREADY(s_axi_control_RREADY),
    .RDATA(s_axi_control_RDATA),
    .RRESP(s_axi_control_RRESP),
    .BVALID(s_axi_control_BVALID),
    .BREADY(s_axi_control_BREADY),
    .BRESP(s_axi_control_BRESP),
    .ACLK(ap_clk),
    .ARESET(ap_rst_n_inv),
    .ACLK_EN(1'b1),
    .rmem0(rmem0),
    .rmem1(rmem1),
    .rmem2(rmem2),
    .rmem3(rmem3),
    .rmem4(rmem4),
    .rmem5(rmem5),
    .rmem6(rmem6),
    .rmem7(rmem7),
    .rmem8(rmem8),
    .rmem9(rmem9),
    .rmem10(rmem10),
    .rmem11(rmem11),
    .rmem12(rmem12),
    .rmem13(rmem13),
    .rmem14(rmem14),
    .rmem15(rmem15),
    .rmem16(rmem16),
    .rmem17(rmem17),
    .rmem18(rmem18),
    .rmem19(rmem19),
    .rmem20(rmem20),
    .rmem21(rmem21),
    .rmem22(rmem22),
    .rmem23(rmem23),
    .rmem24(rmem24),
    .rmem25(rmem25),
    .rmem26(rmem26),
    .rmem27(rmem27),
    .n(n),
    .ap_start(ap_start),
    .interrupt(interrupt),
    .ap_ready(ap_ready),
    .ap_done(ap_done),
    .ap_idle(ap_idle)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qr0_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qr0_vadd_bw__dout),
    .if_empty_n(qr0_vadd_bw__empty_n),
    .if_read(qr0_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qr0_vadd_bw__din),
    .if_full_n(qr0_vadd_bw__full_n),
    .if_write(qr0_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qr10_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qr10_vadd_bw__dout),
    .if_empty_n(qr10_vadd_bw__empty_n),
    .if_read(qr10_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qr10_vadd_bw__din),
    .if_full_n(qr10_vadd_bw__full_n),
    .if_write(qr10_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qr11_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qr11_vadd_bw__dout),
    .if_empty_n(qr11_vadd_bw__empty_n),
    .if_read(qr11_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qr11_vadd_bw__din),
    .if_full_n(qr11_vadd_bw__full_n),
    .if_write(qr11_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qr12_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qr12_vadd_bw__dout),
    .if_empty_n(qr12_vadd_bw__empty_n),
    .if_read(qr12_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qr12_vadd_bw__din),
    .if_full_n(qr12_vadd_bw__full_n),
    .if_write(qr12_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qr13_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qr13_vadd_bw__dout),
    .if_empty_n(qr13_vadd_bw__empty_n),
    .if_read(qr13_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qr13_vadd_bw__din),
    .if_full_n(qr13_vadd_bw__full_n),
    .if_write(qr13_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qr14_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qr14_vadd_bw__dout),
    .if_empty_n(qr14_vadd_bw__empty_n),
    .if_read(qr14_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qr14_vadd_bw__din),
    .if_full_n(qr14_vadd_bw__full_n),
    .if_write(qr14_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qr15_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qr15_vadd_bw__dout),
    .if_empty_n(qr15_vadd_bw__empty_n),
    .if_read(qr15_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qr15_vadd_bw__din),
    .if_full_n(qr15_vadd_bw__full_n),
    .if_write(qr15_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qr16_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qr16_vadd_bw__dout),
    .if_empty_n(qr16_vadd_bw__empty_n),
    .if_read(qr16_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qr16_vadd_bw__din),
    .if_full_n(qr16_vadd_bw__full_n),
    .if_write(qr16_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qr17_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qr17_vadd_bw__dout),
    .if_empty_n(qr17_vadd_bw__empty_n),
    .if_read(qr17_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qr17_vadd_bw__din),
    .if_full_n(qr17_vadd_bw__full_n),
    .if_write(qr17_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qr18_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qr18_vadd_bw__dout),
    .if_empty_n(qr18_vadd_bw__empty_n),
    .if_read(qr18_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qr18_vadd_bw__din),
    .if_full_n(qr18_vadd_bw__full_n),
    .if_write(qr18_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qr19_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qr19_vadd_bw__dout),
    .if_empty_n(qr19_vadd_bw__empty_n),
    .if_read(qr19_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qr19_vadd_bw__din),
    .if_full_n(qr19_vadd_bw__full_n),
    .if_write(qr19_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qr1_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qr1_vadd_bw__dout),
    .if_empty_n(qr1_vadd_bw__empty_n),
    .if_read(qr1_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qr1_vadd_bw__din),
    .if_full_n(qr1_vadd_bw__full_n),
    .if_write(qr1_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qr20_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qr20_vadd_bw__dout),
    .if_empty_n(qr20_vadd_bw__empty_n),
    .if_read(qr20_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qr20_vadd_bw__din),
    .if_full_n(qr20_vadd_bw__full_n),
    .if_write(qr20_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qr21_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qr21_vadd_bw__dout),
    .if_empty_n(qr21_vadd_bw__empty_n),
    .if_read(qr21_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qr21_vadd_bw__din),
    .if_full_n(qr21_vadd_bw__full_n),
    .if_write(qr21_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qr22_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qr22_vadd_bw__dout),
    .if_empty_n(qr22_vadd_bw__empty_n),
    .if_read(qr22_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qr22_vadd_bw__din),
    .if_full_n(qr22_vadd_bw__full_n),
    .if_write(qr22_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qr23_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qr23_vadd_bw__dout),
    .if_empty_n(qr23_vadd_bw__empty_n),
    .if_read(qr23_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qr23_vadd_bw__din),
    .if_full_n(qr23_vadd_bw__full_n),
    .if_write(qr23_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qr24_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qr24_vadd_bw__dout),
    .if_empty_n(qr24_vadd_bw__empty_n),
    .if_read(qr24_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qr24_vadd_bw__din),
    .if_full_n(qr24_vadd_bw__full_n),
    .if_write(qr24_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qr25_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qr25_vadd_bw__dout),
    .if_empty_n(qr25_vadd_bw__empty_n),
    .if_read(qr25_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qr25_vadd_bw__din),
    .if_full_n(qr25_vadd_bw__full_n),
    .if_write(qr25_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qr26_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qr26_vadd_bw__dout),
    .if_empty_n(qr26_vadd_bw__empty_n),
    .if_read(qr26_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qr26_vadd_bw__din),
    .if_full_n(qr26_vadd_bw__full_n),
    .if_write(qr26_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qr27_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qr27_vadd_bw__dout),
    .if_empty_n(qr27_vadd_bw__empty_n),
    .if_read(qr27_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qr27_vadd_bw__din),
    .if_full_n(qr27_vadd_bw__full_n),
    .if_write(qr27_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qr2_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qr2_vadd_bw__dout),
    .if_empty_n(qr2_vadd_bw__empty_n),
    .if_read(qr2_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qr2_vadd_bw__din),
    .if_full_n(qr2_vadd_bw__full_n),
    .if_write(qr2_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qr3_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qr3_vadd_bw__dout),
    .if_empty_n(qr3_vadd_bw__empty_n),
    .if_read(qr3_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qr3_vadd_bw__din),
    .if_full_n(qr3_vadd_bw__full_n),
    .if_write(qr3_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qr4_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qr4_vadd_bw__dout),
    .if_empty_n(qr4_vadd_bw__empty_n),
    .if_read(qr4_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qr4_vadd_bw__din),
    .if_full_n(qr4_vadd_bw__full_n),
    .if_write(qr4_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qr5_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qr5_vadd_bw__dout),
    .if_empty_n(qr5_vadd_bw__empty_n),
    .if_read(qr5_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qr5_vadd_bw__din),
    .if_full_n(qr5_vadd_bw__full_n),
    .if_write(qr5_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qr6_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qr6_vadd_bw__dout),
    .if_empty_n(qr6_vadd_bw__empty_n),
    .if_read(qr6_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qr6_vadd_bw__din),
    .if_full_n(qr6_vadd_bw__full_n),
    .if_write(qr6_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qr7_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qr7_vadd_bw__dout),
    .if_empty_n(qr7_vadd_bw__empty_n),
    .if_read(qr7_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qr7_vadd_bw__din),
    .if_full_n(qr7_vadd_bw__full_n),
    .if_write(qr7_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qr8_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qr8_vadd_bw__dout),
    .if_empty_n(qr8_vadd_bw__empty_n),
    .if_read(qr8_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qr8_vadd_bw__din),
    .if_full_n(qr8_vadd_bw__full_n),
    .if_write(qr8_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qr9_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qr9_vadd_bw__dout),
    .if_empty_n(qr9_vadd_bw__empty_n),
    .if_read(qr9_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qr9_vadd_bw__din),
    .if_full_n(qr9_vadd_bw__full_n),
    .if_write(qr9_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qw0_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qw0_vadd_bw__dout),
    .if_empty_n(qw0_vadd_bw__empty_n),
    .if_read(qw0_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qw0_vadd_bw__din),
    .if_full_n(qw0_vadd_bw__full_n),
    .if_write(qw0_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qw10_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qw10_vadd_bw__dout),
    .if_empty_n(qw10_vadd_bw__empty_n),
    .if_read(qw10_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qw10_vadd_bw__din),
    .if_full_n(qw10_vadd_bw__full_n),
    .if_write(qw10_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qw11_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qw11_vadd_bw__dout),
    .if_empty_n(qw11_vadd_bw__empty_n),
    .if_read(qw11_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qw11_vadd_bw__din),
    .if_full_n(qw11_vadd_bw__full_n),
    .if_write(qw11_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qw12_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qw12_vadd_bw__dout),
    .if_empty_n(qw12_vadd_bw__empty_n),
    .if_read(qw12_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qw12_vadd_bw__din),
    .if_full_n(qw12_vadd_bw__full_n),
    .if_write(qw12_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qw13_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qw13_vadd_bw__dout),
    .if_empty_n(qw13_vadd_bw__empty_n),
    .if_read(qw13_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qw13_vadd_bw__din),
    .if_full_n(qw13_vadd_bw__full_n),
    .if_write(qw13_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qw14_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qw14_vadd_bw__dout),
    .if_empty_n(qw14_vadd_bw__empty_n),
    .if_read(qw14_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qw14_vadd_bw__din),
    .if_full_n(qw14_vadd_bw__full_n),
    .if_write(qw14_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qw15_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qw15_vadd_bw__dout),
    .if_empty_n(qw15_vadd_bw__empty_n),
    .if_read(qw15_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qw15_vadd_bw__din),
    .if_full_n(qw15_vadd_bw__full_n),
    .if_write(qw15_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qw16_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qw16_vadd_bw__dout),
    .if_empty_n(qw16_vadd_bw__empty_n),
    .if_read(qw16_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qw16_vadd_bw__din),
    .if_full_n(qw16_vadd_bw__full_n),
    .if_write(qw16_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qw17_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qw17_vadd_bw__dout),
    .if_empty_n(qw17_vadd_bw__empty_n),
    .if_read(qw17_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qw17_vadd_bw__din),
    .if_full_n(qw17_vadd_bw__full_n),
    .if_write(qw17_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qw18_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qw18_vadd_bw__dout),
    .if_empty_n(qw18_vadd_bw__empty_n),
    .if_read(qw18_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qw18_vadd_bw__din),
    .if_full_n(qw18_vadd_bw__full_n),
    .if_write(qw18_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qw19_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qw19_vadd_bw__dout),
    .if_empty_n(qw19_vadd_bw__empty_n),
    .if_read(qw19_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qw19_vadd_bw__din),
    .if_full_n(qw19_vadd_bw__full_n),
    .if_write(qw19_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qw1_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qw1_vadd_bw__dout),
    .if_empty_n(qw1_vadd_bw__empty_n),
    .if_read(qw1_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qw1_vadd_bw__din),
    .if_full_n(qw1_vadd_bw__full_n),
    .if_write(qw1_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qw20_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qw20_vadd_bw__dout),
    .if_empty_n(qw20_vadd_bw__empty_n),
    .if_read(qw20_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qw20_vadd_bw__din),
    .if_full_n(qw20_vadd_bw__full_n),
    .if_write(qw20_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qw21_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qw21_vadd_bw__dout),
    .if_empty_n(qw21_vadd_bw__empty_n),
    .if_read(qw21_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qw21_vadd_bw__din),
    .if_full_n(qw21_vadd_bw__full_n),
    .if_write(qw21_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qw22_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qw22_vadd_bw__dout),
    .if_empty_n(qw22_vadd_bw__empty_n),
    .if_read(qw22_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qw22_vadd_bw__din),
    .if_full_n(qw22_vadd_bw__full_n),
    .if_write(qw22_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qw23_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qw23_vadd_bw__dout),
    .if_empty_n(qw23_vadd_bw__empty_n),
    .if_read(qw23_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qw23_vadd_bw__din),
    .if_full_n(qw23_vadd_bw__full_n),
    .if_write(qw23_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qw24_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qw24_vadd_bw__dout),
    .if_empty_n(qw24_vadd_bw__empty_n),
    .if_read(qw24_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qw24_vadd_bw__din),
    .if_full_n(qw24_vadd_bw__full_n),
    .if_write(qw24_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qw25_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qw25_vadd_bw__dout),
    .if_empty_n(qw25_vadd_bw__empty_n),
    .if_read(qw25_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qw25_vadd_bw__din),
    .if_full_n(qw25_vadd_bw__full_n),
    .if_write(qw25_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qw26_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qw26_vadd_bw__dout),
    .if_empty_n(qw26_vadd_bw__empty_n),
    .if_read(qw26_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qw26_vadd_bw__din),
    .if_full_n(qw26_vadd_bw__full_n),
    .if_write(qw26_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qw27_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qw27_vadd_bw__dout),
    .if_empty_n(qw27_vadd_bw__empty_n),
    .if_read(qw27_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qw27_vadd_bw__din),
    .if_full_n(qw27_vadd_bw__full_n),
    .if_write(qw27_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qw2_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qw2_vadd_bw__dout),
    .if_empty_n(qw2_vadd_bw__empty_n),
    .if_read(qw2_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qw2_vadd_bw__din),
    .if_full_n(qw2_vadd_bw__full_n),
    .if_write(qw2_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qw3_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qw3_vadd_bw__dout),
    .if_empty_n(qw3_vadd_bw__empty_n),
    .if_read(qw3_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qw3_vadd_bw__din),
    .if_full_n(qw3_vadd_bw__full_n),
    .if_write(qw3_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qw4_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qw4_vadd_bw__dout),
    .if_empty_n(qw4_vadd_bw__empty_n),
    .if_read(qw4_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qw4_vadd_bw__din),
    .if_full_n(qw4_vadd_bw__full_n),
    .if_write(qw4_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qw5_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qw5_vadd_bw__dout),
    .if_empty_n(qw5_vadd_bw__empty_n),
    .if_read(qw5_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qw5_vadd_bw__din),
    .if_full_n(qw5_vadd_bw__full_n),
    .if_write(qw5_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qw6_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qw6_vadd_bw__dout),
    .if_empty_n(qw6_vadd_bw__empty_n),
    .if_read(qw6_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qw6_vadd_bw__din),
    .if_full_n(qw6_vadd_bw__full_n),
    .if_write(qw6_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qw7_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qw7_vadd_bw__dout),
    .if_empty_n(qw7_vadd_bw__empty_n),
    .if_read(qw7_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qw7_vadd_bw__din),
    .if_full_n(qw7_vadd_bw__full_n),
    .if_write(qw7_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qw8_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qw8_vadd_bw__dout),
    .if_empty_n(qw8_vadd_bw__empty_n),
    .if_read(qw8_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qw8_vadd_bw__din),
    .if_full_n(qw8_vadd_bw__full_n),
    .if_write(qw8_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  qw9_vadd_bw
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(qw9_vadd_bw__dout),
    .if_empty_n(qw9_vadd_bw__empty_n),
    .if_read(qw9_vadd_bw__read),
    .if_read_ce(1'b1),
    .if_din(qw9_vadd_bw__din),
    .if_full_n(qw9_vadd_bw__full_n),
    .if_write(qw9_vadd_bw__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) axi_crossbar_2x1
  #(
    .DATA_WIDTH(512),
    .ADDR_WIDTH(64),
    .S_ID_WIDTH(1),
    .M_ID_WIDTH(2),
    .M00_ADDR_WIDTH(64),
    .M00_ISSUE(16),
    .S00_THREADS(1),
    .S01_THREADS(1)
  )
  axi_crossbar_2x1__rmem0
  (
    .clk(ap_clk),
    .rst(ap_rst_n_inv),
    .m00_axi_araddr(m_axi_rmem0_ARADDR),
    .m00_axi_arburst(m_axi_rmem0_ARBURST),
    .m00_axi_arcache(m_axi_rmem0_ARCACHE),
    .m00_axi_arid(m_axi_rmem0_ARID),
    .m00_axi_arlen(m_axi_rmem0_ARLEN),
    .m00_axi_arlock(m_axi_rmem0_ARLOCK),
    .m00_axi_arprot(m_axi_rmem0_ARPROT),
    .m00_axi_arqos(m_axi_rmem0_ARQOS),
    .m00_axi_arready(m_axi_rmem0_ARREADY),
    .m00_axi_arsize(m_axi_rmem0_ARSIZE),
    .m00_axi_arvalid(m_axi_rmem0_ARVALID),
    .m00_axi_awaddr(m_axi_rmem0_AWADDR),
    .m00_axi_awburst(m_axi_rmem0_AWBURST),
    .m00_axi_awcache(m_axi_rmem0_AWCACHE),
    .m00_axi_awid(m_axi_rmem0_AWID),
    .m00_axi_awlen(m_axi_rmem0_AWLEN),
    .m00_axi_awlock(m_axi_rmem0_AWLOCK),
    .m00_axi_awprot(m_axi_rmem0_AWPROT),
    .m00_axi_awqos(m_axi_rmem0_AWQOS),
    .m00_axi_awready(m_axi_rmem0_AWREADY),
    .m00_axi_awsize(m_axi_rmem0_AWSIZE),
    .m00_axi_awvalid(m_axi_rmem0_AWVALID),
    .m00_axi_bid(m_axi_rmem0_BID),
    .m00_axi_bready(m_axi_rmem0_BREADY),
    .m00_axi_bresp(m_axi_rmem0_BRESP),
    .m00_axi_bvalid(m_axi_rmem0_BVALID),
    .m00_axi_rdata(m_axi_rmem0_RDATA),
    .m00_axi_rid(m_axi_rmem0_RID),
    .m00_axi_rlast(m_axi_rmem0_RLAST),
    .m00_axi_rready(m_axi_rmem0_RREADY),
    .m00_axi_rresp(m_axi_rmem0_RRESP),
    .m00_axi_rvalid(m_axi_rmem0_RVALID),
    .m00_axi_wdata(m_axi_rmem0_WDATA),
    .m00_axi_wlast(m_axi_rmem0_WLAST),
    .m00_axi_wready(m_axi_rmem0_WREADY),
    .m00_axi_wstrb(m_axi_rmem0_WSTRB),
    .m00_axi_wvalid(m_axi_rmem0_WVALID),
    .s00_axi_araddr(m_axi_rmem0___Mmap2Stream_0___mmap_ARADDR),
    .s00_axi_arburst(m_axi_rmem0___Mmap2Stream_0___mmap_ARBURST),
    .s00_axi_arcache(m_axi_rmem0___Mmap2Stream_0___mmap_ARCACHE),
    .s00_axi_arid(m_axi_rmem0___Mmap2Stream_0___mmap_ARID),
    .s00_axi_arlen(m_axi_rmem0___Mmap2Stream_0___mmap_ARLEN),
    .s00_axi_arlock(m_axi_rmem0___Mmap2Stream_0___mmap_ARLOCK),
    .s00_axi_arprot(m_axi_rmem0___Mmap2Stream_0___mmap_ARPROT),
    .s00_axi_arqos(m_axi_rmem0___Mmap2Stream_0___mmap_ARQOS),
    .s00_axi_arready(m_axi_rmem0___Mmap2Stream_0___mmap_ARREADY),
    .s00_axi_arsize(m_axi_rmem0___Mmap2Stream_0___mmap_ARSIZE),
    .s00_axi_arvalid(m_axi_rmem0___Mmap2Stream_0___mmap_ARVALID),
    .s00_axi_awaddr(m_axi_rmem0___Mmap2Stream_0___mmap_AWADDR),
    .s00_axi_awburst(m_axi_rmem0___Mmap2Stream_0___mmap_AWBURST),
    .s00_axi_awcache(m_axi_rmem0___Mmap2Stream_0___mmap_AWCACHE),
    .s00_axi_awid(m_axi_rmem0___Mmap2Stream_0___mmap_AWID),
    .s00_axi_awlen(m_axi_rmem0___Mmap2Stream_0___mmap_AWLEN),
    .s00_axi_awlock(m_axi_rmem0___Mmap2Stream_0___mmap_AWLOCK),
    .s00_axi_awprot(m_axi_rmem0___Mmap2Stream_0___mmap_AWPROT),
    .s00_axi_awqos(m_axi_rmem0___Mmap2Stream_0___mmap_AWQOS),
    .s00_axi_awready(m_axi_rmem0___Mmap2Stream_0___mmap_AWREADY),
    .s00_axi_awsize(m_axi_rmem0___Mmap2Stream_0___mmap_AWSIZE),
    .s00_axi_awvalid(m_axi_rmem0___Mmap2Stream_0___mmap_AWVALID),
    .s00_axi_bid(m_axi_rmem0___Mmap2Stream_0___mmap_BID),
    .s00_axi_bready(m_axi_rmem0___Mmap2Stream_0___mmap_BREADY),
    .s00_axi_bresp(m_axi_rmem0___Mmap2Stream_0___mmap_BRESP),
    .s00_axi_bvalid(m_axi_rmem0___Mmap2Stream_0___mmap_BVALID),
    .s00_axi_rdata(m_axi_rmem0___Mmap2Stream_0___mmap_RDATA),
    .s00_axi_rid(m_axi_rmem0___Mmap2Stream_0___mmap_RID),
    .s00_axi_rlast(m_axi_rmem0___Mmap2Stream_0___mmap_RLAST),
    .s00_axi_rready(m_axi_rmem0___Mmap2Stream_0___mmap_RREADY),
    .s00_axi_rresp(m_axi_rmem0___Mmap2Stream_0___mmap_RRESP),
    .s00_axi_rvalid(m_axi_rmem0___Mmap2Stream_0___mmap_RVALID),
    .s00_axi_wdata(m_axi_rmem0___Mmap2Stream_0___mmap_WDATA),
    .s00_axi_wlast(m_axi_rmem0___Mmap2Stream_0___mmap_WLAST),
    .s00_axi_wready(m_axi_rmem0___Mmap2Stream_0___mmap_WREADY),
    .s00_axi_wstrb(m_axi_rmem0___Mmap2Stream_0___mmap_WSTRB),
    .s00_axi_wvalid(m_axi_rmem0___Mmap2Stream_0___mmap_WVALID),
    .s01_axi_araddr(m_axi_rmem0___Stream2Mmap_0___mmap_ARADDR),
    .s01_axi_arburst(m_axi_rmem0___Stream2Mmap_0___mmap_ARBURST),
    .s01_axi_arcache(m_axi_rmem0___Stream2Mmap_0___mmap_ARCACHE),
    .s01_axi_arid(m_axi_rmem0___Stream2Mmap_0___mmap_ARID),
    .s01_axi_arlen(m_axi_rmem0___Stream2Mmap_0___mmap_ARLEN),
    .s01_axi_arlock(m_axi_rmem0___Stream2Mmap_0___mmap_ARLOCK),
    .s01_axi_arprot(m_axi_rmem0___Stream2Mmap_0___mmap_ARPROT),
    .s01_axi_arqos(m_axi_rmem0___Stream2Mmap_0___mmap_ARQOS),
    .s01_axi_arready(m_axi_rmem0___Stream2Mmap_0___mmap_ARREADY),
    .s01_axi_arsize(m_axi_rmem0___Stream2Mmap_0___mmap_ARSIZE),
    .s01_axi_arvalid(m_axi_rmem0___Stream2Mmap_0___mmap_ARVALID),
    .s01_axi_awaddr(m_axi_rmem0___Stream2Mmap_0___mmap_AWADDR),
    .s01_axi_awburst(m_axi_rmem0___Stream2Mmap_0___mmap_AWBURST),
    .s01_axi_awcache(m_axi_rmem0___Stream2Mmap_0___mmap_AWCACHE),
    .s01_axi_awid(m_axi_rmem0___Stream2Mmap_0___mmap_AWID),
    .s01_axi_awlen(m_axi_rmem0___Stream2Mmap_0___mmap_AWLEN),
    .s01_axi_awlock(m_axi_rmem0___Stream2Mmap_0___mmap_AWLOCK),
    .s01_axi_awprot(m_axi_rmem0___Stream2Mmap_0___mmap_AWPROT),
    .s01_axi_awqos(m_axi_rmem0___Stream2Mmap_0___mmap_AWQOS),
    .s01_axi_awready(m_axi_rmem0___Stream2Mmap_0___mmap_AWREADY),
    .s01_axi_awsize(m_axi_rmem0___Stream2Mmap_0___mmap_AWSIZE),
    .s01_axi_awvalid(m_axi_rmem0___Stream2Mmap_0___mmap_AWVALID),
    .s01_axi_bid(m_axi_rmem0___Stream2Mmap_0___mmap_BID),
    .s01_axi_bready(m_axi_rmem0___Stream2Mmap_0___mmap_BREADY),
    .s01_axi_bresp(m_axi_rmem0___Stream2Mmap_0___mmap_BRESP),
    .s01_axi_bvalid(m_axi_rmem0___Stream2Mmap_0___mmap_BVALID),
    .s01_axi_rdata(m_axi_rmem0___Stream2Mmap_0___mmap_RDATA),
    .s01_axi_rid(m_axi_rmem0___Stream2Mmap_0___mmap_RID),
    .s01_axi_rlast(m_axi_rmem0___Stream2Mmap_0___mmap_RLAST),
    .s01_axi_rready(m_axi_rmem0___Stream2Mmap_0___mmap_RREADY),
    .s01_axi_rresp(m_axi_rmem0___Stream2Mmap_0___mmap_RRESP),
    .s01_axi_rvalid(m_axi_rmem0___Stream2Mmap_0___mmap_RVALID),
    .s01_axi_wdata(m_axi_rmem0___Stream2Mmap_0___mmap_WDATA),
    .s01_axi_wlast(m_axi_rmem0___Stream2Mmap_0___mmap_WLAST),
    .s01_axi_wready(m_axi_rmem0___Stream2Mmap_0___mmap_WREADY),
    .s01_axi_wstrb(m_axi_rmem0___Stream2Mmap_0___mmap_WSTRB),
    .s01_axi_wvalid(m_axi_rmem0___Stream2Mmap_0___mmap_WVALID)
  );


  (* keep_hierarchy = "yes" *) axi_crossbar_2x1
  #(
    .DATA_WIDTH(512),
    .ADDR_WIDTH(64),
    .S_ID_WIDTH(1),
    .M_ID_WIDTH(2),
    .M00_ADDR_WIDTH(64),
    .M00_ISSUE(16),
    .S00_THREADS(1),
    .S01_THREADS(1)
  )
  axi_crossbar_2x1__rmem1
  (
    .clk(ap_clk),
    .rst(ap_rst_n_inv),
    .m00_axi_araddr(m_axi_rmem1_ARADDR),
    .m00_axi_arburst(m_axi_rmem1_ARBURST),
    .m00_axi_arcache(m_axi_rmem1_ARCACHE),
    .m00_axi_arid(m_axi_rmem1_ARID),
    .m00_axi_arlen(m_axi_rmem1_ARLEN),
    .m00_axi_arlock(m_axi_rmem1_ARLOCK),
    .m00_axi_arprot(m_axi_rmem1_ARPROT),
    .m00_axi_arqos(m_axi_rmem1_ARQOS),
    .m00_axi_arready(m_axi_rmem1_ARREADY),
    .m00_axi_arsize(m_axi_rmem1_ARSIZE),
    .m00_axi_arvalid(m_axi_rmem1_ARVALID),
    .m00_axi_awaddr(m_axi_rmem1_AWADDR),
    .m00_axi_awburst(m_axi_rmem1_AWBURST),
    .m00_axi_awcache(m_axi_rmem1_AWCACHE),
    .m00_axi_awid(m_axi_rmem1_AWID),
    .m00_axi_awlen(m_axi_rmem1_AWLEN),
    .m00_axi_awlock(m_axi_rmem1_AWLOCK),
    .m00_axi_awprot(m_axi_rmem1_AWPROT),
    .m00_axi_awqos(m_axi_rmem1_AWQOS),
    .m00_axi_awready(m_axi_rmem1_AWREADY),
    .m00_axi_awsize(m_axi_rmem1_AWSIZE),
    .m00_axi_awvalid(m_axi_rmem1_AWVALID),
    .m00_axi_bid(m_axi_rmem1_BID),
    .m00_axi_bready(m_axi_rmem1_BREADY),
    .m00_axi_bresp(m_axi_rmem1_BRESP),
    .m00_axi_bvalid(m_axi_rmem1_BVALID),
    .m00_axi_rdata(m_axi_rmem1_RDATA),
    .m00_axi_rid(m_axi_rmem1_RID),
    .m00_axi_rlast(m_axi_rmem1_RLAST),
    .m00_axi_rready(m_axi_rmem1_RREADY),
    .m00_axi_rresp(m_axi_rmem1_RRESP),
    .m00_axi_rvalid(m_axi_rmem1_RVALID),
    .m00_axi_wdata(m_axi_rmem1_WDATA),
    .m00_axi_wlast(m_axi_rmem1_WLAST),
    .m00_axi_wready(m_axi_rmem1_WREADY),
    .m00_axi_wstrb(m_axi_rmem1_WSTRB),
    .m00_axi_wvalid(m_axi_rmem1_WVALID),
    .s00_axi_araddr(m_axi_rmem1___Mmap2Stream_1___mmap_ARADDR),
    .s00_axi_arburst(m_axi_rmem1___Mmap2Stream_1___mmap_ARBURST),
    .s00_axi_arcache(m_axi_rmem1___Mmap2Stream_1___mmap_ARCACHE),
    .s00_axi_arid(m_axi_rmem1___Mmap2Stream_1___mmap_ARID),
    .s00_axi_arlen(m_axi_rmem1___Mmap2Stream_1___mmap_ARLEN),
    .s00_axi_arlock(m_axi_rmem1___Mmap2Stream_1___mmap_ARLOCK),
    .s00_axi_arprot(m_axi_rmem1___Mmap2Stream_1___mmap_ARPROT),
    .s00_axi_arqos(m_axi_rmem1___Mmap2Stream_1___mmap_ARQOS),
    .s00_axi_arready(m_axi_rmem1___Mmap2Stream_1___mmap_ARREADY),
    .s00_axi_arsize(m_axi_rmem1___Mmap2Stream_1___mmap_ARSIZE),
    .s00_axi_arvalid(m_axi_rmem1___Mmap2Stream_1___mmap_ARVALID),
    .s00_axi_awaddr(m_axi_rmem1___Mmap2Stream_1___mmap_AWADDR),
    .s00_axi_awburst(m_axi_rmem1___Mmap2Stream_1___mmap_AWBURST),
    .s00_axi_awcache(m_axi_rmem1___Mmap2Stream_1___mmap_AWCACHE),
    .s00_axi_awid(m_axi_rmem1___Mmap2Stream_1___mmap_AWID),
    .s00_axi_awlen(m_axi_rmem1___Mmap2Stream_1___mmap_AWLEN),
    .s00_axi_awlock(m_axi_rmem1___Mmap2Stream_1___mmap_AWLOCK),
    .s00_axi_awprot(m_axi_rmem1___Mmap2Stream_1___mmap_AWPROT),
    .s00_axi_awqos(m_axi_rmem1___Mmap2Stream_1___mmap_AWQOS),
    .s00_axi_awready(m_axi_rmem1___Mmap2Stream_1___mmap_AWREADY),
    .s00_axi_awsize(m_axi_rmem1___Mmap2Stream_1___mmap_AWSIZE),
    .s00_axi_awvalid(m_axi_rmem1___Mmap2Stream_1___mmap_AWVALID),
    .s00_axi_bid(m_axi_rmem1___Mmap2Stream_1___mmap_BID),
    .s00_axi_bready(m_axi_rmem1___Mmap2Stream_1___mmap_BREADY),
    .s00_axi_bresp(m_axi_rmem1___Mmap2Stream_1___mmap_BRESP),
    .s00_axi_bvalid(m_axi_rmem1___Mmap2Stream_1___mmap_BVALID),
    .s00_axi_rdata(m_axi_rmem1___Mmap2Stream_1___mmap_RDATA),
    .s00_axi_rid(m_axi_rmem1___Mmap2Stream_1___mmap_RID),
    .s00_axi_rlast(m_axi_rmem1___Mmap2Stream_1___mmap_RLAST),
    .s00_axi_rready(m_axi_rmem1___Mmap2Stream_1___mmap_RREADY),
    .s00_axi_rresp(m_axi_rmem1___Mmap2Stream_1___mmap_RRESP),
    .s00_axi_rvalid(m_axi_rmem1___Mmap2Stream_1___mmap_RVALID),
    .s00_axi_wdata(m_axi_rmem1___Mmap2Stream_1___mmap_WDATA),
    .s00_axi_wlast(m_axi_rmem1___Mmap2Stream_1___mmap_WLAST),
    .s00_axi_wready(m_axi_rmem1___Mmap2Stream_1___mmap_WREADY),
    .s00_axi_wstrb(m_axi_rmem1___Mmap2Stream_1___mmap_WSTRB),
    .s00_axi_wvalid(m_axi_rmem1___Mmap2Stream_1___mmap_WVALID),
    .s01_axi_araddr(m_axi_rmem1___Stream2Mmap_1___mmap_ARADDR),
    .s01_axi_arburst(m_axi_rmem1___Stream2Mmap_1___mmap_ARBURST),
    .s01_axi_arcache(m_axi_rmem1___Stream2Mmap_1___mmap_ARCACHE),
    .s01_axi_arid(m_axi_rmem1___Stream2Mmap_1___mmap_ARID),
    .s01_axi_arlen(m_axi_rmem1___Stream2Mmap_1___mmap_ARLEN),
    .s01_axi_arlock(m_axi_rmem1___Stream2Mmap_1___mmap_ARLOCK),
    .s01_axi_arprot(m_axi_rmem1___Stream2Mmap_1___mmap_ARPROT),
    .s01_axi_arqos(m_axi_rmem1___Stream2Mmap_1___mmap_ARQOS),
    .s01_axi_arready(m_axi_rmem1___Stream2Mmap_1___mmap_ARREADY),
    .s01_axi_arsize(m_axi_rmem1___Stream2Mmap_1___mmap_ARSIZE),
    .s01_axi_arvalid(m_axi_rmem1___Stream2Mmap_1___mmap_ARVALID),
    .s01_axi_awaddr(m_axi_rmem1___Stream2Mmap_1___mmap_AWADDR),
    .s01_axi_awburst(m_axi_rmem1___Stream2Mmap_1___mmap_AWBURST),
    .s01_axi_awcache(m_axi_rmem1___Stream2Mmap_1___mmap_AWCACHE),
    .s01_axi_awid(m_axi_rmem1___Stream2Mmap_1___mmap_AWID),
    .s01_axi_awlen(m_axi_rmem1___Stream2Mmap_1___mmap_AWLEN),
    .s01_axi_awlock(m_axi_rmem1___Stream2Mmap_1___mmap_AWLOCK),
    .s01_axi_awprot(m_axi_rmem1___Stream2Mmap_1___mmap_AWPROT),
    .s01_axi_awqos(m_axi_rmem1___Stream2Mmap_1___mmap_AWQOS),
    .s01_axi_awready(m_axi_rmem1___Stream2Mmap_1___mmap_AWREADY),
    .s01_axi_awsize(m_axi_rmem1___Stream2Mmap_1___mmap_AWSIZE),
    .s01_axi_awvalid(m_axi_rmem1___Stream2Mmap_1___mmap_AWVALID),
    .s01_axi_bid(m_axi_rmem1___Stream2Mmap_1___mmap_BID),
    .s01_axi_bready(m_axi_rmem1___Stream2Mmap_1___mmap_BREADY),
    .s01_axi_bresp(m_axi_rmem1___Stream2Mmap_1___mmap_BRESP),
    .s01_axi_bvalid(m_axi_rmem1___Stream2Mmap_1___mmap_BVALID),
    .s01_axi_rdata(m_axi_rmem1___Stream2Mmap_1___mmap_RDATA),
    .s01_axi_rid(m_axi_rmem1___Stream2Mmap_1___mmap_RID),
    .s01_axi_rlast(m_axi_rmem1___Stream2Mmap_1___mmap_RLAST),
    .s01_axi_rready(m_axi_rmem1___Stream2Mmap_1___mmap_RREADY),
    .s01_axi_rresp(m_axi_rmem1___Stream2Mmap_1___mmap_RRESP),
    .s01_axi_rvalid(m_axi_rmem1___Stream2Mmap_1___mmap_RVALID),
    .s01_axi_wdata(m_axi_rmem1___Stream2Mmap_1___mmap_WDATA),
    .s01_axi_wlast(m_axi_rmem1___Stream2Mmap_1___mmap_WLAST),
    .s01_axi_wready(m_axi_rmem1___Stream2Mmap_1___mmap_WREADY),
    .s01_axi_wstrb(m_axi_rmem1___Stream2Mmap_1___mmap_WSTRB),
    .s01_axi_wvalid(m_axi_rmem1___Stream2Mmap_1___mmap_WVALID)
  );


  (* keep_hierarchy = "yes" *) axi_crossbar_2x1
  #(
    .DATA_WIDTH(512),
    .ADDR_WIDTH(64),
    .S_ID_WIDTH(1),
    .M_ID_WIDTH(2),
    .M00_ADDR_WIDTH(64),
    .M00_ISSUE(16),
    .S00_THREADS(1),
    .S01_THREADS(1)
  )
  axi_crossbar_2x1__rmem2
  (
    .clk(ap_clk),
    .rst(ap_rst_n_inv),
    .m00_axi_araddr(m_axi_rmem2_ARADDR),
    .m00_axi_arburst(m_axi_rmem2_ARBURST),
    .m00_axi_arcache(m_axi_rmem2_ARCACHE),
    .m00_axi_arid(m_axi_rmem2_ARID),
    .m00_axi_arlen(m_axi_rmem2_ARLEN),
    .m00_axi_arlock(m_axi_rmem2_ARLOCK),
    .m00_axi_arprot(m_axi_rmem2_ARPROT),
    .m00_axi_arqos(m_axi_rmem2_ARQOS),
    .m00_axi_arready(m_axi_rmem2_ARREADY),
    .m00_axi_arsize(m_axi_rmem2_ARSIZE),
    .m00_axi_arvalid(m_axi_rmem2_ARVALID),
    .m00_axi_awaddr(m_axi_rmem2_AWADDR),
    .m00_axi_awburst(m_axi_rmem2_AWBURST),
    .m00_axi_awcache(m_axi_rmem2_AWCACHE),
    .m00_axi_awid(m_axi_rmem2_AWID),
    .m00_axi_awlen(m_axi_rmem2_AWLEN),
    .m00_axi_awlock(m_axi_rmem2_AWLOCK),
    .m00_axi_awprot(m_axi_rmem2_AWPROT),
    .m00_axi_awqos(m_axi_rmem2_AWQOS),
    .m00_axi_awready(m_axi_rmem2_AWREADY),
    .m00_axi_awsize(m_axi_rmem2_AWSIZE),
    .m00_axi_awvalid(m_axi_rmem2_AWVALID),
    .m00_axi_bid(m_axi_rmem2_BID),
    .m00_axi_bready(m_axi_rmem2_BREADY),
    .m00_axi_bresp(m_axi_rmem2_BRESP),
    .m00_axi_bvalid(m_axi_rmem2_BVALID),
    .m00_axi_rdata(m_axi_rmem2_RDATA),
    .m00_axi_rid(m_axi_rmem2_RID),
    .m00_axi_rlast(m_axi_rmem2_RLAST),
    .m00_axi_rready(m_axi_rmem2_RREADY),
    .m00_axi_rresp(m_axi_rmem2_RRESP),
    .m00_axi_rvalid(m_axi_rmem2_RVALID),
    .m00_axi_wdata(m_axi_rmem2_WDATA),
    .m00_axi_wlast(m_axi_rmem2_WLAST),
    .m00_axi_wready(m_axi_rmem2_WREADY),
    .m00_axi_wstrb(m_axi_rmem2_WSTRB),
    .m00_axi_wvalid(m_axi_rmem2_WVALID),
    .s00_axi_araddr(m_axi_rmem2___Mmap2Stream_2___mmap_ARADDR),
    .s00_axi_arburst(m_axi_rmem2___Mmap2Stream_2___mmap_ARBURST),
    .s00_axi_arcache(m_axi_rmem2___Mmap2Stream_2___mmap_ARCACHE),
    .s00_axi_arid(m_axi_rmem2___Mmap2Stream_2___mmap_ARID),
    .s00_axi_arlen(m_axi_rmem2___Mmap2Stream_2___mmap_ARLEN),
    .s00_axi_arlock(m_axi_rmem2___Mmap2Stream_2___mmap_ARLOCK),
    .s00_axi_arprot(m_axi_rmem2___Mmap2Stream_2___mmap_ARPROT),
    .s00_axi_arqos(m_axi_rmem2___Mmap2Stream_2___mmap_ARQOS),
    .s00_axi_arready(m_axi_rmem2___Mmap2Stream_2___mmap_ARREADY),
    .s00_axi_arsize(m_axi_rmem2___Mmap2Stream_2___mmap_ARSIZE),
    .s00_axi_arvalid(m_axi_rmem2___Mmap2Stream_2___mmap_ARVALID),
    .s00_axi_awaddr(m_axi_rmem2___Mmap2Stream_2___mmap_AWADDR),
    .s00_axi_awburst(m_axi_rmem2___Mmap2Stream_2___mmap_AWBURST),
    .s00_axi_awcache(m_axi_rmem2___Mmap2Stream_2___mmap_AWCACHE),
    .s00_axi_awid(m_axi_rmem2___Mmap2Stream_2___mmap_AWID),
    .s00_axi_awlen(m_axi_rmem2___Mmap2Stream_2___mmap_AWLEN),
    .s00_axi_awlock(m_axi_rmem2___Mmap2Stream_2___mmap_AWLOCK),
    .s00_axi_awprot(m_axi_rmem2___Mmap2Stream_2___mmap_AWPROT),
    .s00_axi_awqos(m_axi_rmem2___Mmap2Stream_2___mmap_AWQOS),
    .s00_axi_awready(m_axi_rmem2___Mmap2Stream_2___mmap_AWREADY),
    .s00_axi_awsize(m_axi_rmem2___Mmap2Stream_2___mmap_AWSIZE),
    .s00_axi_awvalid(m_axi_rmem2___Mmap2Stream_2___mmap_AWVALID),
    .s00_axi_bid(m_axi_rmem2___Mmap2Stream_2___mmap_BID),
    .s00_axi_bready(m_axi_rmem2___Mmap2Stream_2___mmap_BREADY),
    .s00_axi_bresp(m_axi_rmem2___Mmap2Stream_2___mmap_BRESP),
    .s00_axi_bvalid(m_axi_rmem2___Mmap2Stream_2___mmap_BVALID),
    .s00_axi_rdata(m_axi_rmem2___Mmap2Stream_2___mmap_RDATA),
    .s00_axi_rid(m_axi_rmem2___Mmap2Stream_2___mmap_RID),
    .s00_axi_rlast(m_axi_rmem2___Mmap2Stream_2___mmap_RLAST),
    .s00_axi_rready(m_axi_rmem2___Mmap2Stream_2___mmap_RREADY),
    .s00_axi_rresp(m_axi_rmem2___Mmap2Stream_2___mmap_RRESP),
    .s00_axi_rvalid(m_axi_rmem2___Mmap2Stream_2___mmap_RVALID),
    .s00_axi_wdata(m_axi_rmem2___Mmap2Stream_2___mmap_WDATA),
    .s00_axi_wlast(m_axi_rmem2___Mmap2Stream_2___mmap_WLAST),
    .s00_axi_wready(m_axi_rmem2___Mmap2Stream_2___mmap_WREADY),
    .s00_axi_wstrb(m_axi_rmem2___Mmap2Stream_2___mmap_WSTRB),
    .s00_axi_wvalid(m_axi_rmem2___Mmap2Stream_2___mmap_WVALID),
    .s01_axi_araddr(m_axi_rmem2___Stream2Mmap_2___mmap_ARADDR),
    .s01_axi_arburst(m_axi_rmem2___Stream2Mmap_2___mmap_ARBURST),
    .s01_axi_arcache(m_axi_rmem2___Stream2Mmap_2___mmap_ARCACHE),
    .s01_axi_arid(m_axi_rmem2___Stream2Mmap_2___mmap_ARID),
    .s01_axi_arlen(m_axi_rmem2___Stream2Mmap_2___mmap_ARLEN),
    .s01_axi_arlock(m_axi_rmem2___Stream2Mmap_2___mmap_ARLOCK),
    .s01_axi_arprot(m_axi_rmem2___Stream2Mmap_2___mmap_ARPROT),
    .s01_axi_arqos(m_axi_rmem2___Stream2Mmap_2___mmap_ARQOS),
    .s01_axi_arready(m_axi_rmem2___Stream2Mmap_2___mmap_ARREADY),
    .s01_axi_arsize(m_axi_rmem2___Stream2Mmap_2___mmap_ARSIZE),
    .s01_axi_arvalid(m_axi_rmem2___Stream2Mmap_2___mmap_ARVALID),
    .s01_axi_awaddr(m_axi_rmem2___Stream2Mmap_2___mmap_AWADDR),
    .s01_axi_awburst(m_axi_rmem2___Stream2Mmap_2___mmap_AWBURST),
    .s01_axi_awcache(m_axi_rmem2___Stream2Mmap_2___mmap_AWCACHE),
    .s01_axi_awid(m_axi_rmem2___Stream2Mmap_2___mmap_AWID),
    .s01_axi_awlen(m_axi_rmem2___Stream2Mmap_2___mmap_AWLEN),
    .s01_axi_awlock(m_axi_rmem2___Stream2Mmap_2___mmap_AWLOCK),
    .s01_axi_awprot(m_axi_rmem2___Stream2Mmap_2___mmap_AWPROT),
    .s01_axi_awqos(m_axi_rmem2___Stream2Mmap_2___mmap_AWQOS),
    .s01_axi_awready(m_axi_rmem2___Stream2Mmap_2___mmap_AWREADY),
    .s01_axi_awsize(m_axi_rmem2___Stream2Mmap_2___mmap_AWSIZE),
    .s01_axi_awvalid(m_axi_rmem2___Stream2Mmap_2___mmap_AWVALID),
    .s01_axi_bid(m_axi_rmem2___Stream2Mmap_2___mmap_BID),
    .s01_axi_bready(m_axi_rmem2___Stream2Mmap_2___mmap_BREADY),
    .s01_axi_bresp(m_axi_rmem2___Stream2Mmap_2___mmap_BRESP),
    .s01_axi_bvalid(m_axi_rmem2___Stream2Mmap_2___mmap_BVALID),
    .s01_axi_rdata(m_axi_rmem2___Stream2Mmap_2___mmap_RDATA),
    .s01_axi_rid(m_axi_rmem2___Stream2Mmap_2___mmap_RID),
    .s01_axi_rlast(m_axi_rmem2___Stream2Mmap_2___mmap_RLAST),
    .s01_axi_rready(m_axi_rmem2___Stream2Mmap_2___mmap_RREADY),
    .s01_axi_rresp(m_axi_rmem2___Stream2Mmap_2___mmap_RRESP),
    .s01_axi_rvalid(m_axi_rmem2___Stream2Mmap_2___mmap_RVALID),
    .s01_axi_wdata(m_axi_rmem2___Stream2Mmap_2___mmap_WDATA),
    .s01_axi_wlast(m_axi_rmem2___Stream2Mmap_2___mmap_WLAST),
    .s01_axi_wready(m_axi_rmem2___Stream2Mmap_2___mmap_WREADY),
    .s01_axi_wstrb(m_axi_rmem2___Stream2Mmap_2___mmap_WSTRB),
    .s01_axi_wvalid(m_axi_rmem2___Stream2Mmap_2___mmap_WVALID)
  );


  (* keep_hierarchy = "yes" *) axi_crossbar_2x1
  #(
    .DATA_WIDTH(512),
    .ADDR_WIDTH(64),
    .S_ID_WIDTH(1),
    .M_ID_WIDTH(2),
    .M00_ADDR_WIDTH(64),
    .M00_ISSUE(16),
    .S00_THREADS(1),
    .S01_THREADS(1)
  )
  axi_crossbar_2x1__rmem3
  (
    .clk(ap_clk),
    .rst(ap_rst_n_inv),
    .m00_axi_araddr(m_axi_rmem3_ARADDR),
    .m00_axi_arburst(m_axi_rmem3_ARBURST),
    .m00_axi_arcache(m_axi_rmem3_ARCACHE),
    .m00_axi_arid(m_axi_rmem3_ARID),
    .m00_axi_arlen(m_axi_rmem3_ARLEN),
    .m00_axi_arlock(m_axi_rmem3_ARLOCK),
    .m00_axi_arprot(m_axi_rmem3_ARPROT),
    .m00_axi_arqos(m_axi_rmem3_ARQOS),
    .m00_axi_arready(m_axi_rmem3_ARREADY),
    .m00_axi_arsize(m_axi_rmem3_ARSIZE),
    .m00_axi_arvalid(m_axi_rmem3_ARVALID),
    .m00_axi_awaddr(m_axi_rmem3_AWADDR),
    .m00_axi_awburst(m_axi_rmem3_AWBURST),
    .m00_axi_awcache(m_axi_rmem3_AWCACHE),
    .m00_axi_awid(m_axi_rmem3_AWID),
    .m00_axi_awlen(m_axi_rmem3_AWLEN),
    .m00_axi_awlock(m_axi_rmem3_AWLOCK),
    .m00_axi_awprot(m_axi_rmem3_AWPROT),
    .m00_axi_awqos(m_axi_rmem3_AWQOS),
    .m00_axi_awready(m_axi_rmem3_AWREADY),
    .m00_axi_awsize(m_axi_rmem3_AWSIZE),
    .m00_axi_awvalid(m_axi_rmem3_AWVALID),
    .m00_axi_bid(m_axi_rmem3_BID),
    .m00_axi_bready(m_axi_rmem3_BREADY),
    .m00_axi_bresp(m_axi_rmem3_BRESP),
    .m00_axi_bvalid(m_axi_rmem3_BVALID),
    .m00_axi_rdata(m_axi_rmem3_RDATA),
    .m00_axi_rid(m_axi_rmem3_RID),
    .m00_axi_rlast(m_axi_rmem3_RLAST),
    .m00_axi_rready(m_axi_rmem3_RREADY),
    .m00_axi_rresp(m_axi_rmem3_RRESP),
    .m00_axi_rvalid(m_axi_rmem3_RVALID),
    .m00_axi_wdata(m_axi_rmem3_WDATA),
    .m00_axi_wlast(m_axi_rmem3_WLAST),
    .m00_axi_wready(m_axi_rmem3_WREADY),
    .m00_axi_wstrb(m_axi_rmem3_WSTRB),
    .m00_axi_wvalid(m_axi_rmem3_WVALID),
    .s00_axi_araddr(m_axi_rmem3___Mmap2Stream_3___mmap_ARADDR),
    .s00_axi_arburst(m_axi_rmem3___Mmap2Stream_3___mmap_ARBURST),
    .s00_axi_arcache(m_axi_rmem3___Mmap2Stream_3___mmap_ARCACHE),
    .s00_axi_arid(m_axi_rmem3___Mmap2Stream_3___mmap_ARID),
    .s00_axi_arlen(m_axi_rmem3___Mmap2Stream_3___mmap_ARLEN),
    .s00_axi_arlock(m_axi_rmem3___Mmap2Stream_3___mmap_ARLOCK),
    .s00_axi_arprot(m_axi_rmem3___Mmap2Stream_3___mmap_ARPROT),
    .s00_axi_arqos(m_axi_rmem3___Mmap2Stream_3___mmap_ARQOS),
    .s00_axi_arready(m_axi_rmem3___Mmap2Stream_3___mmap_ARREADY),
    .s00_axi_arsize(m_axi_rmem3___Mmap2Stream_3___mmap_ARSIZE),
    .s00_axi_arvalid(m_axi_rmem3___Mmap2Stream_3___mmap_ARVALID),
    .s00_axi_awaddr(m_axi_rmem3___Mmap2Stream_3___mmap_AWADDR),
    .s00_axi_awburst(m_axi_rmem3___Mmap2Stream_3___mmap_AWBURST),
    .s00_axi_awcache(m_axi_rmem3___Mmap2Stream_3___mmap_AWCACHE),
    .s00_axi_awid(m_axi_rmem3___Mmap2Stream_3___mmap_AWID),
    .s00_axi_awlen(m_axi_rmem3___Mmap2Stream_3___mmap_AWLEN),
    .s00_axi_awlock(m_axi_rmem3___Mmap2Stream_3___mmap_AWLOCK),
    .s00_axi_awprot(m_axi_rmem3___Mmap2Stream_3___mmap_AWPROT),
    .s00_axi_awqos(m_axi_rmem3___Mmap2Stream_3___mmap_AWQOS),
    .s00_axi_awready(m_axi_rmem3___Mmap2Stream_3___mmap_AWREADY),
    .s00_axi_awsize(m_axi_rmem3___Mmap2Stream_3___mmap_AWSIZE),
    .s00_axi_awvalid(m_axi_rmem3___Mmap2Stream_3___mmap_AWVALID),
    .s00_axi_bid(m_axi_rmem3___Mmap2Stream_3___mmap_BID),
    .s00_axi_bready(m_axi_rmem3___Mmap2Stream_3___mmap_BREADY),
    .s00_axi_bresp(m_axi_rmem3___Mmap2Stream_3___mmap_BRESP),
    .s00_axi_bvalid(m_axi_rmem3___Mmap2Stream_3___mmap_BVALID),
    .s00_axi_rdata(m_axi_rmem3___Mmap2Stream_3___mmap_RDATA),
    .s00_axi_rid(m_axi_rmem3___Mmap2Stream_3___mmap_RID),
    .s00_axi_rlast(m_axi_rmem3___Mmap2Stream_3___mmap_RLAST),
    .s00_axi_rready(m_axi_rmem3___Mmap2Stream_3___mmap_RREADY),
    .s00_axi_rresp(m_axi_rmem3___Mmap2Stream_3___mmap_RRESP),
    .s00_axi_rvalid(m_axi_rmem3___Mmap2Stream_3___mmap_RVALID),
    .s00_axi_wdata(m_axi_rmem3___Mmap2Stream_3___mmap_WDATA),
    .s00_axi_wlast(m_axi_rmem3___Mmap2Stream_3___mmap_WLAST),
    .s00_axi_wready(m_axi_rmem3___Mmap2Stream_3___mmap_WREADY),
    .s00_axi_wstrb(m_axi_rmem3___Mmap2Stream_3___mmap_WSTRB),
    .s00_axi_wvalid(m_axi_rmem3___Mmap2Stream_3___mmap_WVALID),
    .s01_axi_araddr(m_axi_rmem3___Stream2Mmap_3___mmap_ARADDR),
    .s01_axi_arburst(m_axi_rmem3___Stream2Mmap_3___mmap_ARBURST),
    .s01_axi_arcache(m_axi_rmem3___Stream2Mmap_3___mmap_ARCACHE),
    .s01_axi_arid(m_axi_rmem3___Stream2Mmap_3___mmap_ARID),
    .s01_axi_arlen(m_axi_rmem3___Stream2Mmap_3___mmap_ARLEN),
    .s01_axi_arlock(m_axi_rmem3___Stream2Mmap_3___mmap_ARLOCK),
    .s01_axi_arprot(m_axi_rmem3___Stream2Mmap_3___mmap_ARPROT),
    .s01_axi_arqos(m_axi_rmem3___Stream2Mmap_3___mmap_ARQOS),
    .s01_axi_arready(m_axi_rmem3___Stream2Mmap_3___mmap_ARREADY),
    .s01_axi_arsize(m_axi_rmem3___Stream2Mmap_3___mmap_ARSIZE),
    .s01_axi_arvalid(m_axi_rmem3___Stream2Mmap_3___mmap_ARVALID),
    .s01_axi_awaddr(m_axi_rmem3___Stream2Mmap_3___mmap_AWADDR),
    .s01_axi_awburst(m_axi_rmem3___Stream2Mmap_3___mmap_AWBURST),
    .s01_axi_awcache(m_axi_rmem3___Stream2Mmap_3___mmap_AWCACHE),
    .s01_axi_awid(m_axi_rmem3___Stream2Mmap_3___mmap_AWID),
    .s01_axi_awlen(m_axi_rmem3___Stream2Mmap_3___mmap_AWLEN),
    .s01_axi_awlock(m_axi_rmem3___Stream2Mmap_3___mmap_AWLOCK),
    .s01_axi_awprot(m_axi_rmem3___Stream2Mmap_3___mmap_AWPROT),
    .s01_axi_awqos(m_axi_rmem3___Stream2Mmap_3___mmap_AWQOS),
    .s01_axi_awready(m_axi_rmem3___Stream2Mmap_3___mmap_AWREADY),
    .s01_axi_awsize(m_axi_rmem3___Stream2Mmap_3___mmap_AWSIZE),
    .s01_axi_awvalid(m_axi_rmem3___Stream2Mmap_3___mmap_AWVALID),
    .s01_axi_bid(m_axi_rmem3___Stream2Mmap_3___mmap_BID),
    .s01_axi_bready(m_axi_rmem3___Stream2Mmap_3___mmap_BREADY),
    .s01_axi_bresp(m_axi_rmem3___Stream2Mmap_3___mmap_BRESP),
    .s01_axi_bvalid(m_axi_rmem3___Stream2Mmap_3___mmap_BVALID),
    .s01_axi_rdata(m_axi_rmem3___Stream2Mmap_3___mmap_RDATA),
    .s01_axi_rid(m_axi_rmem3___Stream2Mmap_3___mmap_RID),
    .s01_axi_rlast(m_axi_rmem3___Stream2Mmap_3___mmap_RLAST),
    .s01_axi_rready(m_axi_rmem3___Stream2Mmap_3___mmap_RREADY),
    .s01_axi_rresp(m_axi_rmem3___Stream2Mmap_3___mmap_RRESP),
    .s01_axi_rvalid(m_axi_rmem3___Stream2Mmap_3___mmap_RVALID),
    .s01_axi_wdata(m_axi_rmem3___Stream2Mmap_3___mmap_WDATA),
    .s01_axi_wlast(m_axi_rmem3___Stream2Mmap_3___mmap_WLAST),
    .s01_axi_wready(m_axi_rmem3___Stream2Mmap_3___mmap_WREADY),
    .s01_axi_wstrb(m_axi_rmem3___Stream2Mmap_3___mmap_WSTRB),
    .s01_axi_wvalid(m_axi_rmem3___Stream2Mmap_3___mmap_WVALID)
  );


  (* keep_hierarchy = "yes" *) axi_crossbar_2x1
  #(
    .DATA_WIDTH(512),
    .ADDR_WIDTH(64),
    .S_ID_WIDTH(1),
    .M_ID_WIDTH(2),
    .M00_ADDR_WIDTH(64),
    .M00_ISSUE(16),
    .S00_THREADS(1),
    .S01_THREADS(1)
  )
  axi_crossbar_2x1__rmem4
  (
    .clk(ap_clk),
    .rst(ap_rst_n_inv),
    .m00_axi_araddr(m_axi_rmem4_ARADDR),
    .m00_axi_arburst(m_axi_rmem4_ARBURST),
    .m00_axi_arcache(m_axi_rmem4_ARCACHE),
    .m00_axi_arid(m_axi_rmem4_ARID),
    .m00_axi_arlen(m_axi_rmem4_ARLEN),
    .m00_axi_arlock(m_axi_rmem4_ARLOCK),
    .m00_axi_arprot(m_axi_rmem4_ARPROT),
    .m00_axi_arqos(m_axi_rmem4_ARQOS),
    .m00_axi_arready(m_axi_rmem4_ARREADY),
    .m00_axi_arsize(m_axi_rmem4_ARSIZE),
    .m00_axi_arvalid(m_axi_rmem4_ARVALID),
    .m00_axi_awaddr(m_axi_rmem4_AWADDR),
    .m00_axi_awburst(m_axi_rmem4_AWBURST),
    .m00_axi_awcache(m_axi_rmem4_AWCACHE),
    .m00_axi_awid(m_axi_rmem4_AWID),
    .m00_axi_awlen(m_axi_rmem4_AWLEN),
    .m00_axi_awlock(m_axi_rmem4_AWLOCK),
    .m00_axi_awprot(m_axi_rmem4_AWPROT),
    .m00_axi_awqos(m_axi_rmem4_AWQOS),
    .m00_axi_awready(m_axi_rmem4_AWREADY),
    .m00_axi_awsize(m_axi_rmem4_AWSIZE),
    .m00_axi_awvalid(m_axi_rmem4_AWVALID),
    .m00_axi_bid(m_axi_rmem4_BID),
    .m00_axi_bready(m_axi_rmem4_BREADY),
    .m00_axi_bresp(m_axi_rmem4_BRESP),
    .m00_axi_bvalid(m_axi_rmem4_BVALID),
    .m00_axi_rdata(m_axi_rmem4_RDATA),
    .m00_axi_rid(m_axi_rmem4_RID),
    .m00_axi_rlast(m_axi_rmem4_RLAST),
    .m00_axi_rready(m_axi_rmem4_RREADY),
    .m00_axi_rresp(m_axi_rmem4_RRESP),
    .m00_axi_rvalid(m_axi_rmem4_RVALID),
    .m00_axi_wdata(m_axi_rmem4_WDATA),
    .m00_axi_wlast(m_axi_rmem4_WLAST),
    .m00_axi_wready(m_axi_rmem4_WREADY),
    .m00_axi_wstrb(m_axi_rmem4_WSTRB),
    .m00_axi_wvalid(m_axi_rmem4_WVALID),
    .s00_axi_araddr(m_axi_rmem4___Mmap2Stream_4___mmap_ARADDR),
    .s00_axi_arburst(m_axi_rmem4___Mmap2Stream_4___mmap_ARBURST),
    .s00_axi_arcache(m_axi_rmem4___Mmap2Stream_4___mmap_ARCACHE),
    .s00_axi_arid(m_axi_rmem4___Mmap2Stream_4___mmap_ARID),
    .s00_axi_arlen(m_axi_rmem4___Mmap2Stream_4___mmap_ARLEN),
    .s00_axi_arlock(m_axi_rmem4___Mmap2Stream_4___mmap_ARLOCK),
    .s00_axi_arprot(m_axi_rmem4___Mmap2Stream_4___mmap_ARPROT),
    .s00_axi_arqos(m_axi_rmem4___Mmap2Stream_4___mmap_ARQOS),
    .s00_axi_arready(m_axi_rmem4___Mmap2Stream_4___mmap_ARREADY),
    .s00_axi_arsize(m_axi_rmem4___Mmap2Stream_4___mmap_ARSIZE),
    .s00_axi_arvalid(m_axi_rmem4___Mmap2Stream_4___mmap_ARVALID),
    .s00_axi_awaddr(m_axi_rmem4___Mmap2Stream_4___mmap_AWADDR),
    .s00_axi_awburst(m_axi_rmem4___Mmap2Stream_4___mmap_AWBURST),
    .s00_axi_awcache(m_axi_rmem4___Mmap2Stream_4___mmap_AWCACHE),
    .s00_axi_awid(m_axi_rmem4___Mmap2Stream_4___mmap_AWID),
    .s00_axi_awlen(m_axi_rmem4___Mmap2Stream_4___mmap_AWLEN),
    .s00_axi_awlock(m_axi_rmem4___Mmap2Stream_4___mmap_AWLOCK),
    .s00_axi_awprot(m_axi_rmem4___Mmap2Stream_4___mmap_AWPROT),
    .s00_axi_awqos(m_axi_rmem4___Mmap2Stream_4___mmap_AWQOS),
    .s00_axi_awready(m_axi_rmem4___Mmap2Stream_4___mmap_AWREADY),
    .s00_axi_awsize(m_axi_rmem4___Mmap2Stream_4___mmap_AWSIZE),
    .s00_axi_awvalid(m_axi_rmem4___Mmap2Stream_4___mmap_AWVALID),
    .s00_axi_bid(m_axi_rmem4___Mmap2Stream_4___mmap_BID),
    .s00_axi_bready(m_axi_rmem4___Mmap2Stream_4___mmap_BREADY),
    .s00_axi_bresp(m_axi_rmem4___Mmap2Stream_4___mmap_BRESP),
    .s00_axi_bvalid(m_axi_rmem4___Mmap2Stream_4___mmap_BVALID),
    .s00_axi_rdata(m_axi_rmem4___Mmap2Stream_4___mmap_RDATA),
    .s00_axi_rid(m_axi_rmem4___Mmap2Stream_4___mmap_RID),
    .s00_axi_rlast(m_axi_rmem4___Mmap2Stream_4___mmap_RLAST),
    .s00_axi_rready(m_axi_rmem4___Mmap2Stream_4___mmap_RREADY),
    .s00_axi_rresp(m_axi_rmem4___Mmap2Stream_4___mmap_RRESP),
    .s00_axi_rvalid(m_axi_rmem4___Mmap2Stream_4___mmap_RVALID),
    .s00_axi_wdata(m_axi_rmem4___Mmap2Stream_4___mmap_WDATA),
    .s00_axi_wlast(m_axi_rmem4___Mmap2Stream_4___mmap_WLAST),
    .s00_axi_wready(m_axi_rmem4___Mmap2Stream_4___mmap_WREADY),
    .s00_axi_wstrb(m_axi_rmem4___Mmap2Stream_4___mmap_WSTRB),
    .s00_axi_wvalid(m_axi_rmem4___Mmap2Stream_4___mmap_WVALID),
    .s01_axi_araddr(m_axi_rmem4___Stream2Mmap_4___mmap_ARADDR),
    .s01_axi_arburst(m_axi_rmem4___Stream2Mmap_4___mmap_ARBURST),
    .s01_axi_arcache(m_axi_rmem4___Stream2Mmap_4___mmap_ARCACHE),
    .s01_axi_arid(m_axi_rmem4___Stream2Mmap_4___mmap_ARID),
    .s01_axi_arlen(m_axi_rmem4___Stream2Mmap_4___mmap_ARLEN),
    .s01_axi_arlock(m_axi_rmem4___Stream2Mmap_4___mmap_ARLOCK),
    .s01_axi_arprot(m_axi_rmem4___Stream2Mmap_4___mmap_ARPROT),
    .s01_axi_arqos(m_axi_rmem4___Stream2Mmap_4___mmap_ARQOS),
    .s01_axi_arready(m_axi_rmem4___Stream2Mmap_4___mmap_ARREADY),
    .s01_axi_arsize(m_axi_rmem4___Stream2Mmap_4___mmap_ARSIZE),
    .s01_axi_arvalid(m_axi_rmem4___Stream2Mmap_4___mmap_ARVALID),
    .s01_axi_awaddr(m_axi_rmem4___Stream2Mmap_4___mmap_AWADDR),
    .s01_axi_awburst(m_axi_rmem4___Stream2Mmap_4___mmap_AWBURST),
    .s01_axi_awcache(m_axi_rmem4___Stream2Mmap_4___mmap_AWCACHE),
    .s01_axi_awid(m_axi_rmem4___Stream2Mmap_4___mmap_AWID),
    .s01_axi_awlen(m_axi_rmem4___Stream2Mmap_4___mmap_AWLEN),
    .s01_axi_awlock(m_axi_rmem4___Stream2Mmap_4___mmap_AWLOCK),
    .s01_axi_awprot(m_axi_rmem4___Stream2Mmap_4___mmap_AWPROT),
    .s01_axi_awqos(m_axi_rmem4___Stream2Mmap_4___mmap_AWQOS),
    .s01_axi_awready(m_axi_rmem4___Stream2Mmap_4___mmap_AWREADY),
    .s01_axi_awsize(m_axi_rmem4___Stream2Mmap_4___mmap_AWSIZE),
    .s01_axi_awvalid(m_axi_rmem4___Stream2Mmap_4___mmap_AWVALID),
    .s01_axi_bid(m_axi_rmem4___Stream2Mmap_4___mmap_BID),
    .s01_axi_bready(m_axi_rmem4___Stream2Mmap_4___mmap_BREADY),
    .s01_axi_bresp(m_axi_rmem4___Stream2Mmap_4___mmap_BRESP),
    .s01_axi_bvalid(m_axi_rmem4___Stream2Mmap_4___mmap_BVALID),
    .s01_axi_rdata(m_axi_rmem4___Stream2Mmap_4___mmap_RDATA),
    .s01_axi_rid(m_axi_rmem4___Stream2Mmap_4___mmap_RID),
    .s01_axi_rlast(m_axi_rmem4___Stream2Mmap_4___mmap_RLAST),
    .s01_axi_rready(m_axi_rmem4___Stream2Mmap_4___mmap_RREADY),
    .s01_axi_rresp(m_axi_rmem4___Stream2Mmap_4___mmap_RRESP),
    .s01_axi_rvalid(m_axi_rmem4___Stream2Mmap_4___mmap_RVALID),
    .s01_axi_wdata(m_axi_rmem4___Stream2Mmap_4___mmap_WDATA),
    .s01_axi_wlast(m_axi_rmem4___Stream2Mmap_4___mmap_WLAST),
    .s01_axi_wready(m_axi_rmem4___Stream2Mmap_4___mmap_WREADY),
    .s01_axi_wstrb(m_axi_rmem4___Stream2Mmap_4___mmap_WSTRB),
    .s01_axi_wvalid(m_axi_rmem4___Stream2Mmap_4___mmap_WVALID)
  );


  (* keep_hierarchy = "yes" *) axi_crossbar_2x1
  #(
    .DATA_WIDTH(512),
    .ADDR_WIDTH(64),
    .S_ID_WIDTH(1),
    .M_ID_WIDTH(2),
    .M00_ADDR_WIDTH(64),
    .M00_ISSUE(16),
    .S00_THREADS(1),
    .S01_THREADS(1)
  )
  axi_crossbar_2x1__rmem5
  (
    .clk(ap_clk),
    .rst(ap_rst_n_inv),
    .m00_axi_araddr(m_axi_rmem5_ARADDR),
    .m00_axi_arburst(m_axi_rmem5_ARBURST),
    .m00_axi_arcache(m_axi_rmem5_ARCACHE),
    .m00_axi_arid(m_axi_rmem5_ARID),
    .m00_axi_arlen(m_axi_rmem5_ARLEN),
    .m00_axi_arlock(m_axi_rmem5_ARLOCK),
    .m00_axi_arprot(m_axi_rmem5_ARPROT),
    .m00_axi_arqos(m_axi_rmem5_ARQOS),
    .m00_axi_arready(m_axi_rmem5_ARREADY),
    .m00_axi_arsize(m_axi_rmem5_ARSIZE),
    .m00_axi_arvalid(m_axi_rmem5_ARVALID),
    .m00_axi_awaddr(m_axi_rmem5_AWADDR),
    .m00_axi_awburst(m_axi_rmem5_AWBURST),
    .m00_axi_awcache(m_axi_rmem5_AWCACHE),
    .m00_axi_awid(m_axi_rmem5_AWID),
    .m00_axi_awlen(m_axi_rmem5_AWLEN),
    .m00_axi_awlock(m_axi_rmem5_AWLOCK),
    .m00_axi_awprot(m_axi_rmem5_AWPROT),
    .m00_axi_awqos(m_axi_rmem5_AWQOS),
    .m00_axi_awready(m_axi_rmem5_AWREADY),
    .m00_axi_awsize(m_axi_rmem5_AWSIZE),
    .m00_axi_awvalid(m_axi_rmem5_AWVALID),
    .m00_axi_bid(m_axi_rmem5_BID),
    .m00_axi_bready(m_axi_rmem5_BREADY),
    .m00_axi_bresp(m_axi_rmem5_BRESP),
    .m00_axi_bvalid(m_axi_rmem5_BVALID),
    .m00_axi_rdata(m_axi_rmem5_RDATA),
    .m00_axi_rid(m_axi_rmem5_RID),
    .m00_axi_rlast(m_axi_rmem5_RLAST),
    .m00_axi_rready(m_axi_rmem5_RREADY),
    .m00_axi_rresp(m_axi_rmem5_RRESP),
    .m00_axi_rvalid(m_axi_rmem5_RVALID),
    .m00_axi_wdata(m_axi_rmem5_WDATA),
    .m00_axi_wlast(m_axi_rmem5_WLAST),
    .m00_axi_wready(m_axi_rmem5_WREADY),
    .m00_axi_wstrb(m_axi_rmem5_WSTRB),
    .m00_axi_wvalid(m_axi_rmem5_WVALID),
    .s00_axi_araddr(m_axi_rmem5___Mmap2Stream_5___mmap_ARADDR),
    .s00_axi_arburst(m_axi_rmem5___Mmap2Stream_5___mmap_ARBURST),
    .s00_axi_arcache(m_axi_rmem5___Mmap2Stream_5___mmap_ARCACHE),
    .s00_axi_arid(m_axi_rmem5___Mmap2Stream_5___mmap_ARID),
    .s00_axi_arlen(m_axi_rmem5___Mmap2Stream_5___mmap_ARLEN),
    .s00_axi_arlock(m_axi_rmem5___Mmap2Stream_5___mmap_ARLOCK),
    .s00_axi_arprot(m_axi_rmem5___Mmap2Stream_5___mmap_ARPROT),
    .s00_axi_arqos(m_axi_rmem5___Mmap2Stream_5___mmap_ARQOS),
    .s00_axi_arready(m_axi_rmem5___Mmap2Stream_5___mmap_ARREADY),
    .s00_axi_arsize(m_axi_rmem5___Mmap2Stream_5___mmap_ARSIZE),
    .s00_axi_arvalid(m_axi_rmem5___Mmap2Stream_5___mmap_ARVALID),
    .s00_axi_awaddr(m_axi_rmem5___Mmap2Stream_5___mmap_AWADDR),
    .s00_axi_awburst(m_axi_rmem5___Mmap2Stream_5___mmap_AWBURST),
    .s00_axi_awcache(m_axi_rmem5___Mmap2Stream_5___mmap_AWCACHE),
    .s00_axi_awid(m_axi_rmem5___Mmap2Stream_5___mmap_AWID),
    .s00_axi_awlen(m_axi_rmem5___Mmap2Stream_5___mmap_AWLEN),
    .s00_axi_awlock(m_axi_rmem5___Mmap2Stream_5___mmap_AWLOCK),
    .s00_axi_awprot(m_axi_rmem5___Mmap2Stream_5___mmap_AWPROT),
    .s00_axi_awqos(m_axi_rmem5___Mmap2Stream_5___mmap_AWQOS),
    .s00_axi_awready(m_axi_rmem5___Mmap2Stream_5___mmap_AWREADY),
    .s00_axi_awsize(m_axi_rmem5___Mmap2Stream_5___mmap_AWSIZE),
    .s00_axi_awvalid(m_axi_rmem5___Mmap2Stream_5___mmap_AWVALID),
    .s00_axi_bid(m_axi_rmem5___Mmap2Stream_5___mmap_BID),
    .s00_axi_bready(m_axi_rmem5___Mmap2Stream_5___mmap_BREADY),
    .s00_axi_bresp(m_axi_rmem5___Mmap2Stream_5___mmap_BRESP),
    .s00_axi_bvalid(m_axi_rmem5___Mmap2Stream_5___mmap_BVALID),
    .s00_axi_rdata(m_axi_rmem5___Mmap2Stream_5___mmap_RDATA),
    .s00_axi_rid(m_axi_rmem5___Mmap2Stream_5___mmap_RID),
    .s00_axi_rlast(m_axi_rmem5___Mmap2Stream_5___mmap_RLAST),
    .s00_axi_rready(m_axi_rmem5___Mmap2Stream_5___mmap_RREADY),
    .s00_axi_rresp(m_axi_rmem5___Mmap2Stream_5___mmap_RRESP),
    .s00_axi_rvalid(m_axi_rmem5___Mmap2Stream_5___mmap_RVALID),
    .s00_axi_wdata(m_axi_rmem5___Mmap2Stream_5___mmap_WDATA),
    .s00_axi_wlast(m_axi_rmem5___Mmap2Stream_5___mmap_WLAST),
    .s00_axi_wready(m_axi_rmem5___Mmap2Stream_5___mmap_WREADY),
    .s00_axi_wstrb(m_axi_rmem5___Mmap2Stream_5___mmap_WSTRB),
    .s00_axi_wvalid(m_axi_rmem5___Mmap2Stream_5___mmap_WVALID),
    .s01_axi_araddr(m_axi_rmem5___Stream2Mmap_5___mmap_ARADDR),
    .s01_axi_arburst(m_axi_rmem5___Stream2Mmap_5___mmap_ARBURST),
    .s01_axi_arcache(m_axi_rmem5___Stream2Mmap_5___mmap_ARCACHE),
    .s01_axi_arid(m_axi_rmem5___Stream2Mmap_5___mmap_ARID),
    .s01_axi_arlen(m_axi_rmem5___Stream2Mmap_5___mmap_ARLEN),
    .s01_axi_arlock(m_axi_rmem5___Stream2Mmap_5___mmap_ARLOCK),
    .s01_axi_arprot(m_axi_rmem5___Stream2Mmap_5___mmap_ARPROT),
    .s01_axi_arqos(m_axi_rmem5___Stream2Mmap_5___mmap_ARQOS),
    .s01_axi_arready(m_axi_rmem5___Stream2Mmap_5___mmap_ARREADY),
    .s01_axi_arsize(m_axi_rmem5___Stream2Mmap_5___mmap_ARSIZE),
    .s01_axi_arvalid(m_axi_rmem5___Stream2Mmap_5___mmap_ARVALID),
    .s01_axi_awaddr(m_axi_rmem5___Stream2Mmap_5___mmap_AWADDR),
    .s01_axi_awburst(m_axi_rmem5___Stream2Mmap_5___mmap_AWBURST),
    .s01_axi_awcache(m_axi_rmem5___Stream2Mmap_5___mmap_AWCACHE),
    .s01_axi_awid(m_axi_rmem5___Stream2Mmap_5___mmap_AWID),
    .s01_axi_awlen(m_axi_rmem5___Stream2Mmap_5___mmap_AWLEN),
    .s01_axi_awlock(m_axi_rmem5___Stream2Mmap_5___mmap_AWLOCK),
    .s01_axi_awprot(m_axi_rmem5___Stream2Mmap_5___mmap_AWPROT),
    .s01_axi_awqos(m_axi_rmem5___Stream2Mmap_5___mmap_AWQOS),
    .s01_axi_awready(m_axi_rmem5___Stream2Mmap_5___mmap_AWREADY),
    .s01_axi_awsize(m_axi_rmem5___Stream2Mmap_5___mmap_AWSIZE),
    .s01_axi_awvalid(m_axi_rmem5___Stream2Mmap_5___mmap_AWVALID),
    .s01_axi_bid(m_axi_rmem5___Stream2Mmap_5___mmap_BID),
    .s01_axi_bready(m_axi_rmem5___Stream2Mmap_5___mmap_BREADY),
    .s01_axi_bresp(m_axi_rmem5___Stream2Mmap_5___mmap_BRESP),
    .s01_axi_bvalid(m_axi_rmem5___Stream2Mmap_5___mmap_BVALID),
    .s01_axi_rdata(m_axi_rmem5___Stream2Mmap_5___mmap_RDATA),
    .s01_axi_rid(m_axi_rmem5___Stream2Mmap_5___mmap_RID),
    .s01_axi_rlast(m_axi_rmem5___Stream2Mmap_5___mmap_RLAST),
    .s01_axi_rready(m_axi_rmem5___Stream2Mmap_5___mmap_RREADY),
    .s01_axi_rresp(m_axi_rmem5___Stream2Mmap_5___mmap_RRESP),
    .s01_axi_rvalid(m_axi_rmem5___Stream2Mmap_5___mmap_RVALID),
    .s01_axi_wdata(m_axi_rmem5___Stream2Mmap_5___mmap_WDATA),
    .s01_axi_wlast(m_axi_rmem5___Stream2Mmap_5___mmap_WLAST),
    .s01_axi_wready(m_axi_rmem5___Stream2Mmap_5___mmap_WREADY),
    .s01_axi_wstrb(m_axi_rmem5___Stream2Mmap_5___mmap_WSTRB),
    .s01_axi_wvalid(m_axi_rmem5___Stream2Mmap_5___mmap_WVALID)
  );


  (* keep_hierarchy = "yes" *) axi_crossbar_2x1
  #(
    .DATA_WIDTH(512),
    .ADDR_WIDTH(64),
    .S_ID_WIDTH(1),
    .M_ID_WIDTH(2),
    .M00_ADDR_WIDTH(64),
    .M00_ISSUE(16),
    .S00_THREADS(1),
    .S01_THREADS(1)
  )
  axi_crossbar_2x1__rmem6
  (
    .clk(ap_clk),
    .rst(ap_rst_n_inv),
    .m00_axi_araddr(m_axi_rmem6_ARADDR),
    .m00_axi_arburst(m_axi_rmem6_ARBURST),
    .m00_axi_arcache(m_axi_rmem6_ARCACHE),
    .m00_axi_arid(m_axi_rmem6_ARID),
    .m00_axi_arlen(m_axi_rmem6_ARLEN),
    .m00_axi_arlock(m_axi_rmem6_ARLOCK),
    .m00_axi_arprot(m_axi_rmem6_ARPROT),
    .m00_axi_arqos(m_axi_rmem6_ARQOS),
    .m00_axi_arready(m_axi_rmem6_ARREADY),
    .m00_axi_arsize(m_axi_rmem6_ARSIZE),
    .m00_axi_arvalid(m_axi_rmem6_ARVALID),
    .m00_axi_awaddr(m_axi_rmem6_AWADDR),
    .m00_axi_awburst(m_axi_rmem6_AWBURST),
    .m00_axi_awcache(m_axi_rmem6_AWCACHE),
    .m00_axi_awid(m_axi_rmem6_AWID),
    .m00_axi_awlen(m_axi_rmem6_AWLEN),
    .m00_axi_awlock(m_axi_rmem6_AWLOCK),
    .m00_axi_awprot(m_axi_rmem6_AWPROT),
    .m00_axi_awqos(m_axi_rmem6_AWQOS),
    .m00_axi_awready(m_axi_rmem6_AWREADY),
    .m00_axi_awsize(m_axi_rmem6_AWSIZE),
    .m00_axi_awvalid(m_axi_rmem6_AWVALID),
    .m00_axi_bid(m_axi_rmem6_BID),
    .m00_axi_bready(m_axi_rmem6_BREADY),
    .m00_axi_bresp(m_axi_rmem6_BRESP),
    .m00_axi_bvalid(m_axi_rmem6_BVALID),
    .m00_axi_rdata(m_axi_rmem6_RDATA),
    .m00_axi_rid(m_axi_rmem6_RID),
    .m00_axi_rlast(m_axi_rmem6_RLAST),
    .m00_axi_rready(m_axi_rmem6_RREADY),
    .m00_axi_rresp(m_axi_rmem6_RRESP),
    .m00_axi_rvalid(m_axi_rmem6_RVALID),
    .m00_axi_wdata(m_axi_rmem6_WDATA),
    .m00_axi_wlast(m_axi_rmem6_WLAST),
    .m00_axi_wready(m_axi_rmem6_WREADY),
    .m00_axi_wstrb(m_axi_rmem6_WSTRB),
    .m00_axi_wvalid(m_axi_rmem6_WVALID),
    .s00_axi_araddr(m_axi_rmem6___Mmap2Stream_6___mmap_ARADDR),
    .s00_axi_arburst(m_axi_rmem6___Mmap2Stream_6___mmap_ARBURST),
    .s00_axi_arcache(m_axi_rmem6___Mmap2Stream_6___mmap_ARCACHE),
    .s00_axi_arid(m_axi_rmem6___Mmap2Stream_6___mmap_ARID),
    .s00_axi_arlen(m_axi_rmem6___Mmap2Stream_6___mmap_ARLEN),
    .s00_axi_arlock(m_axi_rmem6___Mmap2Stream_6___mmap_ARLOCK),
    .s00_axi_arprot(m_axi_rmem6___Mmap2Stream_6___mmap_ARPROT),
    .s00_axi_arqos(m_axi_rmem6___Mmap2Stream_6___mmap_ARQOS),
    .s00_axi_arready(m_axi_rmem6___Mmap2Stream_6___mmap_ARREADY),
    .s00_axi_arsize(m_axi_rmem6___Mmap2Stream_6___mmap_ARSIZE),
    .s00_axi_arvalid(m_axi_rmem6___Mmap2Stream_6___mmap_ARVALID),
    .s00_axi_awaddr(m_axi_rmem6___Mmap2Stream_6___mmap_AWADDR),
    .s00_axi_awburst(m_axi_rmem6___Mmap2Stream_6___mmap_AWBURST),
    .s00_axi_awcache(m_axi_rmem6___Mmap2Stream_6___mmap_AWCACHE),
    .s00_axi_awid(m_axi_rmem6___Mmap2Stream_6___mmap_AWID),
    .s00_axi_awlen(m_axi_rmem6___Mmap2Stream_6___mmap_AWLEN),
    .s00_axi_awlock(m_axi_rmem6___Mmap2Stream_6___mmap_AWLOCK),
    .s00_axi_awprot(m_axi_rmem6___Mmap2Stream_6___mmap_AWPROT),
    .s00_axi_awqos(m_axi_rmem6___Mmap2Stream_6___mmap_AWQOS),
    .s00_axi_awready(m_axi_rmem6___Mmap2Stream_6___mmap_AWREADY),
    .s00_axi_awsize(m_axi_rmem6___Mmap2Stream_6___mmap_AWSIZE),
    .s00_axi_awvalid(m_axi_rmem6___Mmap2Stream_6___mmap_AWVALID),
    .s00_axi_bid(m_axi_rmem6___Mmap2Stream_6___mmap_BID),
    .s00_axi_bready(m_axi_rmem6___Mmap2Stream_6___mmap_BREADY),
    .s00_axi_bresp(m_axi_rmem6___Mmap2Stream_6___mmap_BRESP),
    .s00_axi_bvalid(m_axi_rmem6___Mmap2Stream_6___mmap_BVALID),
    .s00_axi_rdata(m_axi_rmem6___Mmap2Stream_6___mmap_RDATA),
    .s00_axi_rid(m_axi_rmem6___Mmap2Stream_6___mmap_RID),
    .s00_axi_rlast(m_axi_rmem6___Mmap2Stream_6___mmap_RLAST),
    .s00_axi_rready(m_axi_rmem6___Mmap2Stream_6___mmap_RREADY),
    .s00_axi_rresp(m_axi_rmem6___Mmap2Stream_6___mmap_RRESP),
    .s00_axi_rvalid(m_axi_rmem6___Mmap2Stream_6___mmap_RVALID),
    .s00_axi_wdata(m_axi_rmem6___Mmap2Stream_6___mmap_WDATA),
    .s00_axi_wlast(m_axi_rmem6___Mmap2Stream_6___mmap_WLAST),
    .s00_axi_wready(m_axi_rmem6___Mmap2Stream_6___mmap_WREADY),
    .s00_axi_wstrb(m_axi_rmem6___Mmap2Stream_6___mmap_WSTRB),
    .s00_axi_wvalid(m_axi_rmem6___Mmap2Stream_6___mmap_WVALID),
    .s01_axi_araddr(m_axi_rmem6___Stream2Mmap_6___mmap_ARADDR),
    .s01_axi_arburst(m_axi_rmem6___Stream2Mmap_6___mmap_ARBURST),
    .s01_axi_arcache(m_axi_rmem6___Stream2Mmap_6___mmap_ARCACHE),
    .s01_axi_arid(m_axi_rmem6___Stream2Mmap_6___mmap_ARID),
    .s01_axi_arlen(m_axi_rmem6___Stream2Mmap_6___mmap_ARLEN),
    .s01_axi_arlock(m_axi_rmem6___Stream2Mmap_6___mmap_ARLOCK),
    .s01_axi_arprot(m_axi_rmem6___Stream2Mmap_6___mmap_ARPROT),
    .s01_axi_arqos(m_axi_rmem6___Stream2Mmap_6___mmap_ARQOS),
    .s01_axi_arready(m_axi_rmem6___Stream2Mmap_6___mmap_ARREADY),
    .s01_axi_arsize(m_axi_rmem6___Stream2Mmap_6___mmap_ARSIZE),
    .s01_axi_arvalid(m_axi_rmem6___Stream2Mmap_6___mmap_ARVALID),
    .s01_axi_awaddr(m_axi_rmem6___Stream2Mmap_6___mmap_AWADDR),
    .s01_axi_awburst(m_axi_rmem6___Stream2Mmap_6___mmap_AWBURST),
    .s01_axi_awcache(m_axi_rmem6___Stream2Mmap_6___mmap_AWCACHE),
    .s01_axi_awid(m_axi_rmem6___Stream2Mmap_6___mmap_AWID),
    .s01_axi_awlen(m_axi_rmem6___Stream2Mmap_6___mmap_AWLEN),
    .s01_axi_awlock(m_axi_rmem6___Stream2Mmap_6___mmap_AWLOCK),
    .s01_axi_awprot(m_axi_rmem6___Stream2Mmap_6___mmap_AWPROT),
    .s01_axi_awqos(m_axi_rmem6___Stream2Mmap_6___mmap_AWQOS),
    .s01_axi_awready(m_axi_rmem6___Stream2Mmap_6___mmap_AWREADY),
    .s01_axi_awsize(m_axi_rmem6___Stream2Mmap_6___mmap_AWSIZE),
    .s01_axi_awvalid(m_axi_rmem6___Stream2Mmap_6___mmap_AWVALID),
    .s01_axi_bid(m_axi_rmem6___Stream2Mmap_6___mmap_BID),
    .s01_axi_bready(m_axi_rmem6___Stream2Mmap_6___mmap_BREADY),
    .s01_axi_bresp(m_axi_rmem6___Stream2Mmap_6___mmap_BRESP),
    .s01_axi_bvalid(m_axi_rmem6___Stream2Mmap_6___mmap_BVALID),
    .s01_axi_rdata(m_axi_rmem6___Stream2Mmap_6___mmap_RDATA),
    .s01_axi_rid(m_axi_rmem6___Stream2Mmap_6___mmap_RID),
    .s01_axi_rlast(m_axi_rmem6___Stream2Mmap_6___mmap_RLAST),
    .s01_axi_rready(m_axi_rmem6___Stream2Mmap_6___mmap_RREADY),
    .s01_axi_rresp(m_axi_rmem6___Stream2Mmap_6___mmap_RRESP),
    .s01_axi_rvalid(m_axi_rmem6___Stream2Mmap_6___mmap_RVALID),
    .s01_axi_wdata(m_axi_rmem6___Stream2Mmap_6___mmap_WDATA),
    .s01_axi_wlast(m_axi_rmem6___Stream2Mmap_6___mmap_WLAST),
    .s01_axi_wready(m_axi_rmem6___Stream2Mmap_6___mmap_WREADY),
    .s01_axi_wstrb(m_axi_rmem6___Stream2Mmap_6___mmap_WSTRB),
    .s01_axi_wvalid(m_axi_rmem6___Stream2Mmap_6___mmap_WVALID)
  );


  (* keep_hierarchy = "yes" *) axi_crossbar_2x1
  #(
    .DATA_WIDTH(512),
    .ADDR_WIDTH(64),
    .S_ID_WIDTH(1),
    .M_ID_WIDTH(2),
    .M00_ADDR_WIDTH(64),
    .M00_ISSUE(16),
    .S00_THREADS(1),
    .S01_THREADS(1)
  )
  axi_crossbar_2x1__rmem7
  (
    .clk(ap_clk),
    .rst(ap_rst_n_inv),
    .m00_axi_araddr(m_axi_rmem7_ARADDR),
    .m00_axi_arburst(m_axi_rmem7_ARBURST),
    .m00_axi_arcache(m_axi_rmem7_ARCACHE),
    .m00_axi_arid(m_axi_rmem7_ARID),
    .m00_axi_arlen(m_axi_rmem7_ARLEN),
    .m00_axi_arlock(m_axi_rmem7_ARLOCK),
    .m00_axi_arprot(m_axi_rmem7_ARPROT),
    .m00_axi_arqos(m_axi_rmem7_ARQOS),
    .m00_axi_arready(m_axi_rmem7_ARREADY),
    .m00_axi_arsize(m_axi_rmem7_ARSIZE),
    .m00_axi_arvalid(m_axi_rmem7_ARVALID),
    .m00_axi_awaddr(m_axi_rmem7_AWADDR),
    .m00_axi_awburst(m_axi_rmem7_AWBURST),
    .m00_axi_awcache(m_axi_rmem7_AWCACHE),
    .m00_axi_awid(m_axi_rmem7_AWID),
    .m00_axi_awlen(m_axi_rmem7_AWLEN),
    .m00_axi_awlock(m_axi_rmem7_AWLOCK),
    .m00_axi_awprot(m_axi_rmem7_AWPROT),
    .m00_axi_awqos(m_axi_rmem7_AWQOS),
    .m00_axi_awready(m_axi_rmem7_AWREADY),
    .m00_axi_awsize(m_axi_rmem7_AWSIZE),
    .m00_axi_awvalid(m_axi_rmem7_AWVALID),
    .m00_axi_bid(m_axi_rmem7_BID),
    .m00_axi_bready(m_axi_rmem7_BREADY),
    .m00_axi_bresp(m_axi_rmem7_BRESP),
    .m00_axi_bvalid(m_axi_rmem7_BVALID),
    .m00_axi_rdata(m_axi_rmem7_RDATA),
    .m00_axi_rid(m_axi_rmem7_RID),
    .m00_axi_rlast(m_axi_rmem7_RLAST),
    .m00_axi_rready(m_axi_rmem7_RREADY),
    .m00_axi_rresp(m_axi_rmem7_RRESP),
    .m00_axi_rvalid(m_axi_rmem7_RVALID),
    .m00_axi_wdata(m_axi_rmem7_WDATA),
    .m00_axi_wlast(m_axi_rmem7_WLAST),
    .m00_axi_wready(m_axi_rmem7_WREADY),
    .m00_axi_wstrb(m_axi_rmem7_WSTRB),
    .m00_axi_wvalid(m_axi_rmem7_WVALID),
    .s00_axi_araddr(m_axi_rmem7___Mmap2Stream_7___mmap_ARADDR),
    .s00_axi_arburst(m_axi_rmem7___Mmap2Stream_7___mmap_ARBURST),
    .s00_axi_arcache(m_axi_rmem7___Mmap2Stream_7___mmap_ARCACHE),
    .s00_axi_arid(m_axi_rmem7___Mmap2Stream_7___mmap_ARID),
    .s00_axi_arlen(m_axi_rmem7___Mmap2Stream_7___mmap_ARLEN),
    .s00_axi_arlock(m_axi_rmem7___Mmap2Stream_7___mmap_ARLOCK),
    .s00_axi_arprot(m_axi_rmem7___Mmap2Stream_7___mmap_ARPROT),
    .s00_axi_arqos(m_axi_rmem7___Mmap2Stream_7___mmap_ARQOS),
    .s00_axi_arready(m_axi_rmem7___Mmap2Stream_7___mmap_ARREADY),
    .s00_axi_arsize(m_axi_rmem7___Mmap2Stream_7___mmap_ARSIZE),
    .s00_axi_arvalid(m_axi_rmem7___Mmap2Stream_7___mmap_ARVALID),
    .s00_axi_awaddr(m_axi_rmem7___Mmap2Stream_7___mmap_AWADDR),
    .s00_axi_awburst(m_axi_rmem7___Mmap2Stream_7___mmap_AWBURST),
    .s00_axi_awcache(m_axi_rmem7___Mmap2Stream_7___mmap_AWCACHE),
    .s00_axi_awid(m_axi_rmem7___Mmap2Stream_7___mmap_AWID),
    .s00_axi_awlen(m_axi_rmem7___Mmap2Stream_7___mmap_AWLEN),
    .s00_axi_awlock(m_axi_rmem7___Mmap2Stream_7___mmap_AWLOCK),
    .s00_axi_awprot(m_axi_rmem7___Mmap2Stream_7___mmap_AWPROT),
    .s00_axi_awqos(m_axi_rmem7___Mmap2Stream_7___mmap_AWQOS),
    .s00_axi_awready(m_axi_rmem7___Mmap2Stream_7___mmap_AWREADY),
    .s00_axi_awsize(m_axi_rmem7___Mmap2Stream_7___mmap_AWSIZE),
    .s00_axi_awvalid(m_axi_rmem7___Mmap2Stream_7___mmap_AWVALID),
    .s00_axi_bid(m_axi_rmem7___Mmap2Stream_7___mmap_BID),
    .s00_axi_bready(m_axi_rmem7___Mmap2Stream_7___mmap_BREADY),
    .s00_axi_bresp(m_axi_rmem7___Mmap2Stream_7___mmap_BRESP),
    .s00_axi_bvalid(m_axi_rmem7___Mmap2Stream_7___mmap_BVALID),
    .s00_axi_rdata(m_axi_rmem7___Mmap2Stream_7___mmap_RDATA),
    .s00_axi_rid(m_axi_rmem7___Mmap2Stream_7___mmap_RID),
    .s00_axi_rlast(m_axi_rmem7___Mmap2Stream_7___mmap_RLAST),
    .s00_axi_rready(m_axi_rmem7___Mmap2Stream_7___mmap_RREADY),
    .s00_axi_rresp(m_axi_rmem7___Mmap2Stream_7___mmap_RRESP),
    .s00_axi_rvalid(m_axi_rmem7___Mmap2Stream_7___mmap_RVALID),
    .s00_axi_wdata(m_axi_rmem7___Mmap2Stream_7___mmap_WDATA),
    .s00_axi_wlast(m_axi_rmem7___Mmap2Stream_7___mmap_WLAST),
    .s00_axi_wready(m_axi_rmem7___Mmap2Stream_7___mmap_WREADY),
    .s00_axi_wstrb(m_axi_rmem7___Mmap2Stream_7___mmap_WSTRB),
    .s00_axi_wvalid(m_axi_rmem7___Mmap2Stream_7___mmap_WVALID),
    .s01_axi_araddr(m_axi_rmem7___Stream2Mmap_7___mmap_ARADDR),
    .s01_axi_arburst(m_axi_rmem7___Stream2Mmap_7___mmap_ARBURST),
    .s01_axi_arcache(m_axi_rmem7___Stream2Mmap_7___mmap_ARCACHE),
    .s01_axi_arid(m_axi_rmem7___Stream2Mmap_7___mmap_ARID),
    .s01_axi_arlen(m_axi_rmem7___Stream2Mmap_7___mmap_ARLEN),
    .s01_axi_arlock(m_axi_rmem7___Stream2Mmap_7___mmap_ARLOCK),
    .s01_axi_arprot(m_axi_rmem7___Stream2Mmap_7___mmap_ARPROT),
    .s01_axi_arqos(m_axi_rmem7___Stream2Mmap_7___mmap_ARQOS),
    .s01_axi_arready(m_axi_rmem7___Stream2Mmap_7___mmap_ARREADY),
    .s01_axi_arsize(m_axi_rmem7___Stream2Mmap_7___mmap_ARSIZE),
    .s01_axi_arvalid(m_axi_rmem7___Stream2Mmap_7___mmap_ARVALID),
    .s01_axi_awaddr(m_axi_rmem7___Stream2Mmap_7___mmap_AWADDR),
    .s01_axi_awburst(m_axi_rmem7___Stream2Mmap_7___mmap_AWBURST),
    .s01_axi_awcache(m_axi_rmem7___Stream2Mmap_7___mmap_AWCACHE),
    .s01_axi_awid(m_axi_rmem7___Stream2Mmap_7___mmap_AWID),
    .s01_axi_awlen(m_axi_rmem7___Stream2Mmap_7___mmap_AWLEN),
    .s01_axi_awlock(m_axi_rmem7___Stream2Mmap_7___mmap_AWLOCK),
    .s01_axi_awprot(m_axi_rmem7___Stream2Mmap_7___mmap_AWPROT),
    .s01_axi_awqos(m_axi_rmem7___Stream2Mmap_7___mmap_AWQOS),
    .s01_axi_awready(m_axi_rmem7___Stream2Mmap_7___mmap_AWREADY),
    .s01_axi_awsize(m_axi_rmem7___Stream2Mmap_7___mmap_AWSIZE),
    .s01_axi_awvalid(m_axi_rmem7___Stream2Mmap_7___mmap_AWVALID),
    .s01_axi_bid(m_axi_rmem7___Stream2Mmap_7___mmap_BID),
    .s01_axi_bready(m_axi_rmem7___Stream2Mmap_7___mmap_BREADY),
    .s01_axi_bresp(m_axi_rmem7___Stream2Mmap_7___mmap_BRESP),
    .s01_axi_bvalid(m_axi_rmem7___Stream2Mmap_7___mmap_BVALID),
    .s01_axi_rdata(m_axi_rmem7___Stream2Mmap_7___mmap_RDATA),
    .s01_axi_rid(m_axi_rmem7___Stream2Mmap_7___mmap_RID),
    .s01_axi_rlast(m_axi_rmem7___Stream2Mmap_7___mmap_RLAST),
    .s01_axi_rready(m_axi_rmem7___Stream2Mmap_7___mmap_RREADY),
    .s01_axi_rresp(m_axi_rmem7___Stream2Mmap_7___mmap_RRESP),
    .s01_axi_rvalid(m_axi_rmem7___Stream2Mmap_7___mmap_RVALID),
    .s01_axi_wdata(m_axi_rmem7___Stream2Mmap_7___mmap_WDATA),
    .s01_axi_wlast(m_axi_rmem7___Stream2Mmap_7___mmap_WLAST),
    .s01_axi_wready(m_axi_rmem7___Stream2Mmap_7___mmap_WREADY),
    .s01_axi_wstrb(m_axi_rmem7___Stream2Mmap_7___mmap_WSTRB),
    .s01_axi_wvalid(m_axi_rmem7___Stream2Mmap_7___mmap_WVALID)
  );


  (* keep_hierarchy = "yes" *) axi_crossbar_2x1
  #(
    .DATA_WIDTH(512),
    .ADDR_WIDTH(64),
    .S_ID_WIDTH(1),
    .M_ID_WIDTH(2),
    .M00_ADDR_WIDTH(64),
    .M00_ISSUE(16),
    .S00_THREADS(1),
    .S01_THREADS(1)
  )
  axi_crossbar_2x1__rmem8
  (
    .clk(ap_clk),
    .rst(ap_rst_n_inv),
    .m00_axi_araddr(m_axi_rmem8_ARADDR),
    .m00_axi_arburst(m_axi_rmem8_ARBURST),
    .m00_axi_arcache(m_axi_rmem8_ARCACHE),
    .m00_axi_arid(m_axi_rmem8_ARID),
    .m00_axi_arlen(m_axi_rmem8_ARLEN),
    .m00_axi_arlock(m_axi_rmem8_ARLOCK),
    .m00_axi_arprot(m_axi_rmem8_ARPROT),
    .m00_axi_arqos(m_axi_rmem8_ARQOS),
    .m00_axi_arready(m_axi_rmem8_ARREADY),
    .m00_axi_arsize(m_axi_rmem8_ARSIZE),
    .m00_axi_arvalid(m_axi_rmem8_ARVALID),
    .m00_axi_awaddr(m_axi_rmem8_AWADDR),
    .m00_axi_awburst(m_axi_rmem8_AWBURST),
    .m00_axi_awcache(m_axi_rmem8_AWCACHE),
    .m00_axi_awid(m_axi_rmem8_AWID),
    .m00_axi_awlen(m_axi_rmem8_AWLEN),
    .m00_axi_awlock(m_axi_rmem8_AWLOCK),
    .m00_axi_awprot(m_axi_rmem8_AWPROT),
    .m00_axi_awqos(m_axi_rmem8_AWQOS),
    .m00_axi_awready(m_axi_rmem8_AWREADY),
    .m00_axi_awsize(m_axi_rmem8_AWSIZE),
    .m00_axi_awvalid(m_axi_rmem8_AWVALID),
    .m00_axi_bid(m_axi_rmem8_BID),
    .m00_axi_bready(m_axi_rmem8_BREADY),
    .m00_axi_bresp(m_axi_rmem8_BRESP),
    .m00_axi_bvalid(m_axi_rmem8_BVALID),
    .m00_axi_rdata(m_axi_rmem8_RDATA),
    .m00_axi_rid(m_axi_rmem8_RID),
    .m00_axi_rlast(m_axi_rmem8_RLAST),
    .m00_axi_rready(m_axi_rmem8_RREADY),
    .m00_axi_rresp(m_axi_rmem8_RRESP),
    .m00_axi_rvalid(m_axi_rmem8_RVALID),
    .m00_axi_wdata(m_axi_rmem8_WDATA),
    .m00_axi_wlast(m_axi_rmem8_WLAST),
    .m00_axi_wready(m_axi_rmem8_WREADY),
    .m00_axi_wstrb(m_axi_rmem8_WSTRB),
    .m00_axi_wvalid(m_axi_rmem8_WVALID),
    .s00_axi_araddr(m_axi_rmem8___Mmap2Stream_8___mmap_ARADDR),
    .s00_axi_arburst(m_axi_rmem8___Mmap2Stream_8___mmap_ARBURST),
    .s00_axi_arcache(m_axi_rmem8___Mmap2Stream_8___mmap_ARCACHE),
    .s00_axi_arid(m_axi_rmem8___Mmap2Stream_8___mmap_ARID),
    .s00_axi_arlen(m_axi_rmem8___Mmap2Stream_8___mmap_ARLEN),
    .s00_axi_arlock(m_axi_rmem8___Mmap2Stream_8___mmap_ARLOCK),
    .s00_axi_arprot(m_axi_rmem8___Mmap2Stream_8___mmap_ARPROT),
    .s00_axi_arqos(m_axi_rmem8___Mmap2Stream_8___mmap_ARQOS),
    .s00_axi_arready(m_axi_rmem8___Mmap2Stream_8___mmap_ARREADY),
    .s00_axi_arsize(m_axi_rmem8___Mmap2Stream_8___mmap_ARSIZE),
    .s00_axi_arvalid(m_axi_rmem8___Mmap2Stream_8___mmap_ARVALID),
    .s00_axi_awaddr(m_axi_rmem8___Mmap2Stream_8___mmap_AWADDR),
    .s00_axi_awburst(m_axi_rmem8___Mmap2Stream_8___mmap_AWBURST),
    .s00_axi_awcache(m_axi_rmem8___Mmap2Stream_8___mmap_AWCACHE),
    .s00_axi_awid(m_axi_rmem8___Mmap2Stream_8___mmap_AWID),
    .s00_axi_awlen(m_axi_rmem8___Mmap2Stream_8___mmap_AWLEN),
    .s00_axi_awlock(m_axi_rmem8___Mmap2Stream_8___mmap_AWLOCK),
    .s00_axi_awprot(m_axi_rmem8___Mmap2Stream_8___mmap_AWPROT),
    .s00_axi_awqos(m_axi_rmem8___Mmap2Stream_8___mmap_AWQOS),
    .s00_axi_awready(m_axi_rmem8___Mmap2Stream_8___mmap_AWREADY),
    .s00_axi_awsize(m_axi_rmem8___Mmap2Stream_8___mmap_AWSIZE),
    .s00_axi_awvalid(m_axi_rmem8___Mmap2Stream_8___mmap_AWVALID),
    .s00_axi_bid(m_axi_rmem8___Mmap2Stream_8___mmap_BID),
    .s00_axi_bready(m_axi_rmem8___Mmap2Stream_8___mmap_BREADY),
    .s00_axi_bresp(m_axi_rmem8___Mmap2Stream_8___mmap_BRESP),
    .s00_axi_bvalid(m_axi_rmem8___Mmap2Stream_8___mmap_BVALID),
    .s00_axi_rdata(m_axi_rmem8___Mmap2Stream_8___mmap_RDATA),
    .s00_axi_rid(m_axi_rmem8___Mmap2Stream_8___mmap_RID),
    .s00_axi_rlast(m_axi_rmem8___Mmap2Stream_8___mmap_RLAST),
    .s00_axi_rready(m_axi_rmem8___Mmap2Stream_8___mmap_RREADY),
    .s00_axi_rresp(m_axi_rmem8___Mmap2Stream_8___mmap_RRESP),
    .s00_axi_rvalid(m_axi_rmem8___Mmap2Stream_8___mmap_RVALID),
    .s00_axi_wdata(m_axi_rmem8___Mmap2Stream_8___mmap_WDATA),
    .s00_axi_wlast(m_axi_rmem8___Mmap2Stream_8___mmap_WLAST),
    .s00_axi_wready(m_axi_rmem8___Mmap2Stream_8___mmap_WREADY),
    .s00_axi_wstrb(m_axi_rmem8___Mmap2Stream_8___mmap_WSTRB),
    .s00_axi_wvalid(m_axi_rmem8___Mmap2Stream_8___mmap_WVALID),
    .s01_axi_araddr(m_axi_rmem8___Stream2Mmap_8___mmap_ARADDR),
    .s01_axi_arburst(m_axi_rmem8___Stream2Mmap_8___mmap_ARBURST),
    .s01_axi_arcache(m_axi_rmem8___Stream2Mmap_8___mmap_ARCACHE),
    .s01_axi_arid(m_axi_rmem8___Stream2Mmap_8___mmap_ARID),
    .s01_axi_arlen(m_axi_rmem8___Stream2Mmap_8___mmap_ARLEN),
    .s01_axi_arlock(m_axi_rmem8___Stream2Mmap_8___mmap_ARLOCK),
    .s01_axi_arprot(m_axi_rmem8___Stream2Mmap_8___mmap_ARPROT),
    .s01_axi_arqos(m_axi_rmem8___Stream2Mmap_8___mmap_ARQOS),
    .s01_axi_arready(m_axi_rmem8___Stream2Mmap_8___mmap_ARREADY),
    .s01_axi_arsize(m_axi_rmem8___Stream2Mmap_8___mmap_ARSIZE),
    .s01_axi_arvalid(m_axi_rmem8___Stream2Mmap_8___mmap_ARVALID),
    .s01_axi_awaddr(m_axi_rmem8___Stream2Mmap_8___mmap_AWADDR),
    .s01_axi_awburst(m_axi_rmem8___Stream2Mmap_8___mmap_AWBURST),
    .s01_axi_awcache(m_axi_rmem8___Stream2Mmap_8___mmap_AWCACHE),
    .s01_axi_awid(m_axi_rmem8___Stream2Mmap_8___mmap_AWID),
    .s01_axi_awlen(m_axi_rmem8___Stream2Mmap_8___mmap_AWLEN),
    .s01_axi_awlock(m_axi_rmem8___Stream2Mmap_8___mmap_AWLOCK),
    .s01_axi_awprot(m_axi_rmem8___Stream2Mmap_8___mmap_AWPROT),
    .s01_axi_awqos(m_axi_rmem8___Stream2Mmap_8___mmap_AWQOS),
    .s01_axi_awready(m_axi_rmem8___Stream2Mmap_8___mmap_AWREADY),
    .s01_axi_awsize(m_axi_rmem8___Stream2Mmap_8___mmap_AWSIZE),
    .s01_axi_awvalid(m_axi_rmem8___Stream2Mmap_8___mmap_AWVALID),
    .s01_axi_bid(m_axi_rmem8___Stream2Mmap_8___mmap_BID),
    .s01_axi_bready(m_axi_rmem8___Stream2Mmap_8___mmap_BREADY),
    .s01_axi_bresp(m_axi_rmem8___Stream2Mmap_8___mmap_BRESP),
    .s01_axi_bvalid(m_axi_rmem8___Stream2Mmap_8___mmap_BVALID),
    .s01_axi_rdata(m_axi_rmem8___Stream2Mmap_8___mmap_RDATA),
    .s01_axi_rid(m_axi_rmem8___Stream2Mmap_8___mmap_RID),
    .s01_axi_rlast(m_axi_rmem8___Stream2Mmap_8___mmap_RLAST),
    .s01_axi_rready(m_axi_rmem8___Stream2Mmap_8___mmap_RREADY),
    .s01_axi_rresp(m_axi_rmem8___Stream2Mmap_8___mmap_RRESP),
    .s01_axi_rvalid(m_axi_rmem8___Stream2Mmap_8___mmap_RVALID),
    .s01_axi_wdata(m_axi_rmem8___Stream2Mmap_8___mmap_WDATA),
    .s01_axi_wlast(m_axi_rmem8___Stream2Mmap_8___mmap_WLAST),
    .s01_axi_wready(m_axi_rmem8___Stream2Mmap_8___mmap_WREADY),
    .s01_axi_wstrb(m_axi_rmem8___Stream2Mmap_8___mmap_WSTRB),
    .s01_axi_wvalid(m_axi_rmem8___Stream2Mmap_8___mmap_WVALID)
  );


  (* keep_hierarchy = "yes" *) axi_crossbar_2x1
  #(
    .DATA_WIDTH(512),
    .ADDR_WIDTH(64),
    .S_ID_WIDTH(1),
    .M_ID_WIDTH(2),
    .M00_ADDR_WIDTH(64),
    .M00_ISSUE(16),
    .S00_THREADS(1),
    .S01_THREADS(1)
  )
  axi_crossbar_2x1__rmem9
  (
    .clk(ap_clk),
    .rst(ap_rst_n_inv),
    .m00_axi_araddr(m_axi_rmem9_ARADDR),
    .m00_axi_arburst(m_axi_rmem9_ARBURST),
    .m00_axi_arcache(m_axi_rmem9_ARCACHE),
    .m00_axi_arid(m_axi_rmem9_ARID),
    .m00_axi_arlen(m_axi_rmem9_ARLEN),
    .m00_axi_arlock(m_axi_rmem9_ARLOCK),
    .m00_axi_arprot(m_axi_rmem9_ARPROT),
    .m00_axi_arqos(m_axi_rmem9_ARQOS),
    .m00_axi_arready(m_axi_rmem9_ARREADY),
    .m00_axi_arsize(m_axi_rmem9_ARSIZE),
    .m00_axi_arvalid(m_axi_rmem9_ARVALID),
    .m00_axi_awaddr(m_axi_rmem9_AWADDR),
    .m00_axi_awburst(m_axi_rmem9_AWBURST),
    .m00_axi_awcache(m_axi_rmem9_AWCACHE),
    .m00_axi_awid(m_axi_rmem9_AWID),
    .m00_axi_awlen(m_axi_rmem9_AWLEN),
    .m00_axi_awlock(m_axi_rmem9_AWLOCK),
    .m00_axi_awprot(m_axi_rmem9_AWPROT),
    .m00_axi_awqos(m_axi_rmem9_AWQOS),
    .m00_axi_awready(m_axi_rmem9_AWREADY),
    .m00_axi_awsize(m_axi_rmem9_AWSIZE),
    .m00_axi_awvalid(m_axi_rmem9_AWVALID),
    .m00_axi_bid(m_axi_rmem9_BID),
    .m00_axi_bready(m_axi_rmem9_BREADY),
    .m00_axi_bresp(m_axi_rmem9_BRESP),
    .m00_axi_bvalid(m_axi_rmem9_BVALID),
    .m00_axi_rdata(m_axi_rmem9_RDATA),
    .m00_axi_rid(m_axi_rmem9_RID),
    .m00_axi_rlast(m_axi_rmem9_RLAST),
    .m00_axi_rready(m_axi_rmem9_RREADY),
    .m00_axi_rresp(m_axi_rmem9_RRESP),
    .m00_axi_rvalid(m_axi_rmem9_RVALID),
    .m00_axi_wdata(m_axi_rmem9_WDATA),
    .m00_axi_wlast(m_axi_rmem9_WLAST),
    .m00_axi_wready(m_axi_rmem9_WREADY),
    .m00_axi_wstrb(m_axi_rmem9_WSTRB),
    .m00_axi_wvalid(m_axi_rmem9_WVALID),
    .s00_axi_araddr(m_axi_rmem9___Mmap2Stream_9___mmap_ARADDR),
    .s00_axi_arburst(m_axi_rmem9___Mmap2Stream_9___mmap_ARBURST),
    .s00_axi_arcache(m_axi_rmem9___Mmap2Stream_9___mmap_ARCACHE),
    .s00_axi_arid(m_axi_rmem9___Mmap2Stream_9___mmap_ARID),
    .s00_axi_arlen(m_axi_rmem9___Mmap2Stream_9___mmap_ARLEN),
    .s00_axi_arlock(m_axi_rmem9___Mmap2Stream_9___mmap_ARLOCK),
    .s00_axi_arprot(m_axi_rmem9___Mmap2Stream_9___mmap_ARPROT),
    .s00_axi_arqos(m_axi_rmem9___Mmap2Stream_9___mmap_ARQOS),
    .s00_axi_arready(m_axi_rmem9___Mmap2Stream_9___mmap_ARREADY),
    .s00_axi_arsize(m_axi_rmem9___Mmap2Stream_9___mmap_ARSIZE),
    .s00_axi_arvalid(m_axi_rmem9___Mmap2Stream_9___mmap_ARVALID),
    .s00_axi_awaddr(m_axi_rmem9___Mmap2Stream_9___mmap_AWADDR),
    .s00_axi_awburst(m_axi_rmem9___Mmap2Stream_9___mmap_AWBURST),
    .s00_axi_awcache(m_axi_rmem9___Mmap2Stream_9___mmap_AWCACHE),
    .s00_axi_awid(m_axi_rmem9___Mmap2Stream_9___mmap_AWID),
    .s00_axi_awlen(m_axi_rmem9___Mmap2Stream_9___mmap_AWLEN),
    .s00_axi_awlock(m_axi_rmem9___Mmap2Stream_9___mmap_AWLOCK),
    .s00_axi_awprot(m_axi_rmem9___Mmap2Stream_9___mmap_AWPROT),
    .s00_axi_awqos(m_axi_rmem9___Mmap2Stream_9___mmap_AWQOS),
    .s00_axi_awready(m_axi_rmem9___Mmap2Stream_9___mmap_AWREADY),
    .s00_axi_awsize(m_axi_rmem9___Mmap2Stream_9___mmap_AWSIZE),
    .s00_axi_awvalid(m_axi_rmem9___Mmap2Stream_9___mmap_AWVALID),
    .s00_axi_bid(m_axi_rmem9___Mmap2Stream_9___mmap_BID),
    .s00_axi_bready(m_axi_rmem9___Mmap2Stream_9___mmap_BREADY),
    .s00_axi_bresp(m_axi_rmem9___Mmap2Stream_9___mmap_BRESP),
    .s00_axi_bvalid(m_axi_rmem9___Mmap2Stream_9___mmap_BVALID),
    .s00_axi_rdata(m_axi_rmem9___Mmap2Stream_9___mmap_RDATA),
    .s00_axi_rid(m_axi_rmem9___Mmap2Stream_9___mmap_RID),
    .s00_axi_rlast(m_axi_rmem9___Mmap2Stream_9___mmap_RLAST),
    .s00_axi_rready(m_axi_rmem9___Mmap2Stream_9___mmap_RREADY),
    .s00_axi_rresp(m_axi_rmem9___Mmap2Stream_9___mmap_RRESP),
    .s00_axi_rvalid(m_axi_rmem9___Mmap2Stream_9___mmap_RVALID),
    .s00_axi_wdata(m_axi_rmem9___Mmap2Stream_9___mmap_WDATA),
    .s00_axi_wlast(m_axi_rmem9___Mmap2Stream_9___mmap_WLAST),
    .s00_axi_wready(m_axi_rmem9___Mmap2Stream_9___mmap_WREADY),
    .s00_axi_wstrb(m_axi_rmem9___Mmap2Stream_9___mmap_WSTRB),
    .s00_axi_wvalid(m_axi_rmem9___Mmap2Stream_9___mmap_WVALID),
    .s01_axi_araddr(m_axi_rmem9___Stream2Mmap_9___mmap_ARADDR),
    .s01_axi_arburst(m_axi_rmem9___Stream2Mmap_9___mmap_ARBURST),
    .s01_axi_arcache(m_axi_rmem9___Stream2Mmap_9___mmap_ARCACHE),
    .s01_axi_arid(m_axi_rmem9___Stream2Mmap_9___mmap_ARID),
    .s01_axi_arlen(m_axi_rmem9___Stream2Mmap_9___mmap_ARLEN),
    .s01_axi_arlock(m_axi_rmem9___Stream2Mmap_9___mmap_ARLOCK),
    .s01_axi_arprot(m_axi_rmem9___Stream2Mmap_9___mmap_ARPROT),
    .s01_axi_arqos(m_axi_rmem9___Stream2Mmap_9___mmap_ARQOS),
    .s01_axi_arready(m_axi_rmem9___Stream2Mmap_9___mmap_ARREADY),
    .s01_axi_arsize(m_axi_rmem9___Stream2Mmap_9___mmap_ARSIZE),
    .s01_axi_arvalid(m_axi_rmem9___Stream2Mmap_9___mmap_ARVALID),
    .s01_axi_awaddr(m_axi_rmem9___Stream2Mmap_9___mmap_AWADDR),
    .s01_axi_awburst(m_axi_rmem9___Stream2Mmap_9___mmap_AWBURST),
    .s01_axi_awcache(m_axi_rmem9___Stream2Mmap_9___mmap_AWCACHE),
    .s01_axi_awid(m_axi_rmem9___Stream2Mmap_9___mmap_AWID),
    .s01_axi_awlen(m_axi_rmem9___Stream2Mmap_9___mmap_AWLEN),
    .s01_axi_awlock(m_axi_rmem9___Stream2Mmap_9___mmap_AWLOCK),
    .s01_axi_awprot(m_axi_rmem9___Stream2Mmap_9___mmap_AWPROT),
    .s01_axi_awqos(m_axi_rmem9___Stream2Mmap_9___mmap_AWQOS),
    .s01_axi_awready(m_axi_rmem9___Stream2Mmap_9___mmap_AWREADY),
    .s01_axi_awsize(m_axi_rmem9___Stream2Mmap_9___mmap_AWSIZE),
    .s01_axi_awvalid(m_axi_rmem9___Stream2Mmap_9___mmap_AWVALID),
    .s01_axi_bid(m_axi_rmem9___Stream2Mmap_9___mmap_BID),
    .s01_axi_bready(m_axi_rmem9___Stream2Mmap_9___mmap_BREADY),
    .s01_axi_bresp(m_axi_rmem9___Stream2Mmap_9___mmap_BRESP),
    .s01_axi_bvalid(m_axi_rmem9___Stream2Mmap_9___mmap_BVALID),
    .s01_axi_rdata(m_axi_rmem9___Stream2Mmap_9___mmap_RDATA),
    .s01_axi_rid(m_axi_rmem9___Stream2Mmap_9___mmap_RID),
    .s01_axi_rlast(m_axi_rmem9___Stream2Mmap_9___mmap_RLAST),
    .s01_axi_rready(m_axi_rmem9___Stream2Mmap_9___mmap_RREADY),
    .s01_axi_rresp(m_axi_rmem9___Stream2Mmap_9___mmap_RRESP),
    .s01_axi_rvalid(m_axi_rmem9___Stream2Mmap_9___mmap_RVALID),
    .s01_axi_wdata(m_axi_rmem9___Stream2Mmap_9___mmap_WDATA),
    .s01_axi_wlast(m_axi_rmem9___Stream2Mmap_9___mmap_WLAST),
    .s01_axi_wready(m_axi_rmem9___Stream2Mmap_9___mmap_WREADY),
    .s01_axi_wstrb(m_axi_rmem9___Stream2Mmap_9___mmap_WSTRB),
    .s01_axi_wvalid(m_axi_rmem9___Stream2Mmap_9___mmap_WVALID)
  );


  (* keep_hierarchy = "yes" *) axi_crossbar_2x1
  #(
    .DATA_WIDTH(512),
    .ADDR_WIDTH(64),
    .S_ID_WIDTH(1),
    .M_ID_WIDTH(2),
    .M00_ADDR_WIDTH(64),
    .M00_ISSUE(16),
    .S00_THREADS(1),
    .S01_THREADS(1)
  )
  axi_crossbar_2x1__rmem10
  (
    .clk(ap_clk),
    .rst(ap_rst_n_inv),
    .m00_axi_araddr(m_axi_rmem10_ARADDR),
    .m00_axi_arburst(m_axi_rmem10_ARBURST),
    .m00_axi_arcache(m_axi_rmem10_ARCACHE),
    .m00_axi_arid(m_axi_rmem10_ARID),
    .m00_axi_arlen(m_axi_rmem10_ARLEN),
    .m00_axi_arlock(m_axi_rmem10_ARLOCK),
    .m00_axi_arprot(m_axi_rmem10_ARPROT),
    .m00_axi_arqos(m_axi_rmem10_ARQOS),
    .m00_axi_arready(m_axi_rmem10_ARREADY),
    .m00_axi_arsize(m_axi_rmem10_ARSIZE),
    .m00_axi_arvalid(m_axi_rmem10_ARVALID),
    .m00_axi_awaddr(m_axi_rmem10_AWADDR),
    .m00_axi_awburst(m_axi_rmem10_AWBURST),
    .m00_axi_awcache(m_axi_rmem10_AWCACHE),
    .m00_axi_awid(m_axi_rmem10_AWID),
    .m00_axi_awlen(m_axi_rmem10_AWLEN),
    .m00_axi_awlock(m_axi_rmem10_AWLOCK),
    .m00_axi_awprot(m_axi_rmem10_AWPROT),
    .m00_axi_awqos(m_axi_rmem10_AWQOS),
    .m00_axi_awready(m_axi_rmem10_AWREADY),
    .m00_axi_awsize(m_axi_rmem10_AWSIZE),
    .m00_axi_awvalid(m_axi_rmem10_AWVALID),
    .m00_axi_bid(m_axi_rmem10_BID),
    .m00_axi_bready(m_axi_rmem10_BREADY),
    .m00_axi_bresp(m_axi_rmem10_BRESP),
    .m00_axi_bvalid(m_axi_rmem10_BVALID),
    .m00_axi_rdata(m_axi_rmem10_RDATA),
    .m00_axi_rid(m_axi_rmem10_RID),
    .m00_axi_rlast(m_axi_rmem10_RLAST),
    .m00_axi_rready(m_axi_rmem10_RREADY),
    .m00_axi_rresp(m_axi_rmem10_RRESP),
    .m00_axi_rvalid(m_axi_rmem10_RVALID),
    .m00_axi_wdata(m_axi_rmem10_WDATA),
    .m00_axi_wlast(m_axi_rmem10_WLAST),
    .m00_axi_wready(m_axi_rmem10_WREADY),
    .m00_axi_wstrb(m_axi_rmem10_WSTRB),
    .m00_axi_wvalid(m_axi_rmem10_WVALID),
    .s00_axi_araddr(m_axi_rmem10___Mmap2Stream_10___mmap_ARADDR),
    .s00_axi_arburst(m_axi_rmem10___Mmap2Stream_10___mmap_ARBURST),
    .s00_axi_arcache(m_axi_rmem10___Mmap2Stream_10___mmap_ARCACHE),
    .s00_axi_arid(m_axi_rmem10___Mmap2Stream_10___mmap_ARID),
    .s00_axi_arlen(m_axi_rmem10___Mmap2Stream_10___mmap_ARLEN),
    .s00_axi_arlock(m_axi_rmem10___Mmap2Stream_10___mmap_ARLOCK),
    .s00_axi_arprot(m_axi_rmem10___Mmap2Stream_10___mmap_ARPROT),
    .s00_axi_arqos(m_axi_rmem10___Mmap2Stream_10___mmap_ARQOS),
    .s00_axi_arready(m_axi_rmem10___Mmap2Stream_10___mmap_ARREADY),
    .s00_axi_arsize(m_axi_rmem10___Mmap2Stream_10___mmap_ARSIZE),
    .s00_axi_arvalid(m_axi_rmem10___Mmap2Stream_10___mmap_ARVALID),
    .s00_axi_awaddr(m_axi_rmem10___Mmap2Stream_10___mmap_AWADDR),
    .s00_axi_awburst(m_axi_rmem10___Mmap2Stream_10___mmap_AWBURST),
    .s00_axi_awcache(m_axi_rmem10___Mmap2Stream_10___mmap_AWCACHE),
    .s00_axi_awid(m_axi_rmem10___Mmap2Stream_10___mmap_AWID),
    .s00_axi_awlen(m_axi_rmem10___Mmap2Stream_10___mmap_AWLEN),
    .s00_axi_awlock(m_axi_rmem10___Mmap2Stream_10___mmap_AWLOCK),
    .s00_axi_awprot(m_axi_rmem10___Mmap2Stream_10___mmap_AWPROT),
    .s00_axi_awqos(m_axi_rmem10___Mmap2Stream_10___mmap_AWQOS),
    .s00_axi_awready(m_axi_rmem10___Mmap2Stream_10___mmap_AWREADY),
    .s00_axi_awsize(m_axi_rmem10___Mmap2Stream_10___mmap_AWSIZE),
    .s00_axi_awvalid(m_axi_rmem10___Mmap2Stream_10___mmap_AWVALID),
    .s00_axi_bid(m_axi_rmem10___Mmap2Stream_10___mmap_BID),
    .s00_axi_bready(m_axi_rmem10___Mmap2Stream_10___mmap_BREADY),
    .s00_axi_bresp(m_axi_rmem10___Mmap2Stream_10___mmap_BRESP),
    .s00_axi_bvalid(m_axi_rmem10___Mmap2Stream_10___mmap_BVALID),
    .s00_axi_rdata(m_axi_rmem10___Mmap2Stream_10___mmap_RDATA),
    .s00_axi_rid(m_axi_rmem10___Mmap2Stream_10___mmap_RID),
    .s00_axi_rlast(m_axi_rmem10___Mmap2Stream_10___mmap_RLAST),
    .s00_axi_rready(m_axi_rmem10___Mmap2Stream_10___mmap_RREADY),
    .s00_axi_rresp(m_axi_rmem10___Mmap2Stream_10___mmap_RRESP),
    .s00_axi_rvalid(m_axi_rmem10___Mmap2Stream_10___mmap_RVALID),
    .s00_axi_wdata(m_axi_rmem10___Mmap2Stream_10___mmap_WDATA),
    .s00_axi_wlast(m_axi_rmem10___Mmap2Stream_10___mmap_WLAST),
    .s00_axi_wready(m_axi_rmem10___Mmap2Stream_10___mmap_WREADY),
    .s00_axi_wstrb(m_axi_rmem10___Mmap2Stream_10___mmap_WSTRB),
    .s00_axi_wvalid(m_axi_rmem10___Mmap2Stream_10___mmap_WVALID),
    .s01_axi_araddr(m_axi_rmem10___Stream2Mmap_10___mmap_ARADDR),
    .s01_axi_arburst(m_axi_rmem10___Stream2Mmap_10___mmap_ARBURST),
    .s01_axi_arcache(m_axi_rmem10___Stream2Mmap_10___mmap_ARCACHE),
    .s01_axi_arid(m_axi_rmem10___Stream2Mmap_10___mmap_ARID),
    .s01_axi_arlen(m_axi_rmem10___Stream2Mmap_10___mmap_ARLEN),
    .s01_axi_arlock(m_axi_rmem10___Stream2Mmap_10___mmap_ARLOCK),
    .s01_axi_arprot(m_axi_rmem10___Stream2Mmap_10___mmap_ARPROT),
    .s01_axi_arqos(m_axi_rmem10___Stream2Mmap_10___mmap_ARQOS),
    .s01_axi_arready(m_axi_rmem10___Stream2Mmap_10___mmap_ARREADY),
    .s01_axi_arsize(m_axi_rmem10___Stream2Mmap_10___mmap_ARSIZE),
    .s01_axi_arvalid(m_axi_rmem10___Stream2Mmap_10___mmap_ARVALID),
    .s01_axi_awaddr(m_axi_rmem10___Stream2Mmap_10___mmap_AWADDR),
    .s01_axi_awburst(m_axi_rmem10___Stream2Mmap_10___mmap_AWBURST),
    .s01_axi_awcache(m_axi_rmem10___Stream2Mmap_10___mmap_AWCACHE),
    .s01_axi_awid(m_axi_rmem10___Stream2Mmap_10___mmap_AWID),
    .s01_axi_awlen(m_axi_rmem10___Stream2Mmap_10___mmap_AWLEN),
    .s01_axi_awlock(m_axi_rmem10___Stream2Mmap_10___mmap_AWLOCK),
    .s01_axi_awprot(m_axi_rmem10___Stream2Mmap_10___mmap_AWPROT),
    .s01_axi_awqos(m_axi_rmem10___Stream2Mmap_10___mmap_AWQOS),
    .s01_axi_awready(m_axi_rmem10___Stream2Mmap_10___mmap_AWREADY),
    .s01_axi_awsize(m_axi_rmem10___Stream2Mmap_10___mmap_AWSIZE),
    .s01_axi_awvalid(m_axi_rmem10___Stream2Mmap_10___mmap_AWVALID),
    .s01_axi_bid(m_axi_rmem10___Stream2Mmap_10___mmap_BID),
    .s01_axi_bready(m_axi_rmem10___Stream2Mmap_10___mmap_BREADY),
    .s01_axi_bresp(m_axi_rmem10___Stream2Mmap_10___mmap_BRESP),
    .s01_axi_bvalid(m_axi_rmem10___Stream2Mmap_10___mmap_BVALID),
    .s01_axi_rdata(m_axi_rmem10___Stream2Mmap_10___mmap_RDATA),
    .s01_axi_rid(m_axi_rmem10___Stream2Mmap_10___mmap_RID),
    .s01_axi_rlast(m_axi_rmem10___Stream2Mmap_10___mmap_RLAST),
    .s01_axi_rready(m_axi_rmem10___Stream2Mmap_10___mmap_RREADY),
    .s01_axi_rresp(m_axi_rmem10___Stream2Mmap_10___mmap_RRESP),
    .s01_axi_rvalid(m_axi_rmem10___Stream2Mmap_10___mmap_RVALID),
    .s01_axi_wdata(m_axi_rmem10___Stream2Mmap_10___mmap_WDATA),
    .s01_axi_wlast(m_axi_rmem10___Stream2Mmap_10___mmap_WLAST),
    .s01_axi_wready(m_axi_rmem10___Stream2Mmap_10___mmap_WREADY),
    .s01_axi_wstrb(m_axi_rmem10___Stream2Mmap_10___mmap_WSTRB),
    .s01_axi_wvalid(m_axi_rmem10___Stream2Mmap_10___mmap_WVALID)
  );


  (* keep_hierarchy = "yes" *) axi_crossbar_2x1
  #(
    .DATA_WIDTH(512),
    .ADDR_WIDTH(64),
    .S_ID_WIDTH(1),
    .M_ID_WIDTH(2),
    .M00_ADDR_WIDTH(64),
    .M00_ISSUE(16),
    .S00_THREADS(1),
    .S01_THREADS(1)
  )
  axi_crossbar_2x1__rmem11
  (
    .clk(ap_clk),
    .rst(ap_rst_n_inv),
    .m00_axi_araddr(m_axi_rmem11_ARADDR),
    .m00_axi_arburst(m_axi_rmem11_ARBURST),
    .m00_axi_arcache(m_axi_rmem11_ARCACHE),
    .m00_axi_arid(m_axi_rmem11_ARID),
    .m00_axi_arlen(m_axi_rmem11_ARLEN),
    .m00_axi_arlock(m_axi_rmem11_ARLOCK),
    .m00_axi_arprot(m_axi_rmem11_ARPROT),
    .m00_axi_arqos(m_axi_rmem11_ARQOS),
    .m00_axi_arready(m_axi_rmem11_ARREADY),
    .m00_axi_arsize(m_axi_rmem11_ARSIZE),
    .m00_axi_arvalid(m_axi_rmem11_ARVALID),
    .m00_axi_awaddr(m_axi_rmem11_AWADDR),
    .m00_axi_awburst(m_axi_rmem11_AWBURST),
    .m00_axi_awcache(m_axi_rmem11_AWCACHE),
    .m00_axi_awid(m_axi_rmem11_AWID),
    .m00_axi_awlen(m_axi_rmem11_AWLEN),
    .m00_axi_awlock(m_axi_rmem11_AWLOCK),
    .m00_axi_awprot(m_axi_rmem11_AWPROT),
    .m00_axi_awqos(m_axi_rmem11_AWQOS),
    .m00_axi_awready(m_axi_rmem11_AWREADY),
    .m00_axi_awsize(m_axi_rmem11_AWSIZE),
    .m00_axi_awvalid(m_axi_rmem11_AWVALID),
    .m00_axi_bid(m_axi_rmem11_BID),
    .m00_axi_bready(m_axi_rmem11_BREADY),
    .m00_axi_bresp(m_axi_rmem11_BRESP),
    .m00_axi_bvalid(m_axi_rmem11_BVALID),
    .m00_axi_rdata(m_axi_rmem11_RDATA),
    .m00_axi_rid(m_axi_rmem11_RID),
    .m00_axi_rlast(m_axi_rmem11_RLAST),
    .m00_axi_rready(m_axi_rmem11_RREADY),
    .m00_axi_rresp(m_axi_rmem11_RRESP),
    .m00_axi_rvalid(m_axi_rmem11_RVALID),
    .m00_axi_wdata(m_axi_rmem11_WDATA),
    .m00_axi_wlast(m_axi_rmem11_WLAST),
    .m00_axi_wready(m_axi_rmem11_WREADY),
    .m00_axi_wstrb(m_axi_rmem11_WSTRB),
    .m00_axi_wvalid(m_axi_rmem11_WVALID),
    .s00_axi_araddr(m_axi_rmem11___Mmap2Stream_11___mmap_ARADDR),
    .s00_axi_arburst(m_axi_rmem11___Mmap2Stream_11___mmap_ARBURST),
    .s00_axi_arcache(m_axi_rmem11___Mmap2Stream_11___mmap_ARCACHE),
    .s00_axi_arid(m_axi_rmem11___Mmap2Stream_11___mmap_ARID),
    .s00_axi_arlen(m_axi_rmem11___Mmap2Stream_11___mmap_ARLEN),
    .s00_axi_arlock(m_axi_rmem11___Mmap2Stream_11___mmap_ARLOCK),
    .s00_axi_arprot(m_axi_rmem11___Mmap2Stream_11___mmap_ARPROT),
    .s00_axi_arqos(m_axi_rmem11___Mmap2Stream_11___mmap_ARQOS),
    .s00_axi_arready(m_axi_rmem11___Mmap2Stream_11___mmap_ARREADY),
    .s00_axi_arsize(m_axi_rmem11___Mmap2Stream_11___mmap_ARSIZE),
    .s00_axi_arvalid(m_axi_rmem11___Mmap2Stream_11___mmap_ARVALID),
    .s00_axi_awaddr(m_axi_rmem11___Mmap2Stream_11___mmap_AWADDR),
    .s00_axi_awburst(m_axi_rmem11___Mmap2Stream_11___mmap_AWBURST),
    .s00_axi_awcache(m_axi_rmem11___Mmap2Stream_11___mmap_AWCACHE),
    .s00_axi_awid(m_axi_rmem11___Mmap2Stream_11___mmap_AWID),
    .s00_axi_awlen(m_axi_rmem11___Mmap2Stream_11___mmap_AWLEN),
    .s00_axi_awlock(m_axi_rmem11___Mmap2Stream_11___mmap_AWLOCK),
    .s00_axi_awprot(m_axi_rmem11___Mmap2Stream_11___mmap_AWPROT),
    .s00_axi_awqos(m_axi_rmem11___Mmap2Stream_11___mmap_AWQOS),
    .s00_axi_awready(m_axi_rmem11___Mmap2Stream_11___mmap_AWREADY),
    .s00_axi_awsize(m_axi_rmem11___Mmap2Stream_11___mmap_AWSIZE),
    .s00_axi_awvalid(m_axi_rmem11___Mmap2Stream_11___mmap_AWVALID),
    .s00_axi_bid(m_axi_rmem11___Mmap2Stream_11___mmap_BID),
    .s00_axi_bready(m_axi_rmem11___Mmap2Stream_11___mmap_BREADY),
    .s00_axi_bresp(m_axi_rmem11___Mmap2Stream_11___mmap_BRESP),
    .s00_axi_bvalid(m_axi_rmem11___Mmap2Stream_11___mmap_BVALID),
    .s00_axi_rdata(m_axi_rmem11___Mmap2Stream_11___mmap_RDATA),
    .s00_axi_rid(m_axi_rmem11___Mmap2Stream_11___mmap_RID),
    .s00_axi_rlast(m_axi_rmem11___Mmap2Stream_11___mmap_RLAST),
    .s00_axi_rready(m_axi_rmem11___Mmap2Stream_11___mmap_RREADY),
    .s00_axi_rresp(m_axi_rmem11___Mmap2Stream_11___mmap_RRESP),
    .s00_axi_rvalid(m_axi_rmem11___Mmap2Stream_11___mmap_RVALID),
    .s00_axi_wdata(m_axi_rmem11___Mmap2Stream_11___mmap_WDATA),
    .s00_axi_wlast(m_axi_rmem11___Mmap2Stream_11___mmap_WLAST),
    .s00_axi_wready(m_axi_rmem11___Mmap2Stream_11___mmap_WREADY),
    .s00_axi_wstrb(m_axi_rmem11___Mmap2Stream_11___mmap_WSTRB),
    .s00_axi_wvalid(m_axi_rmem11___Mmap2Stream_11___mmap_WVALID),
    .s01_axi_araddr(m_axi_rmem11___Stream2Mmap_11___mmap_ARADDR),
    .s01_axi_arburst(m_axi_rmem11___Stream2Mmap_11___mmap_ARBURST),
    .s01_axi_arcache(m_axi_rmem11___Stream2Mmap_11___mmap_ARCACHE),
    .s01_axi_arid(m_axi_rmem11___Stream2Mmap_11___mmap_ARID),
    .s01_axi_arlen(m_axi_rmem11___Stream2Mmap_11___mmap_ARLEN),
    .s01_axi_arlock(m_axi_rmem11___Stream2Mmap_11___mmap_ARLOCK),
    .s01_axi_arprot(m_axi_rmem11___Stream2Mmap_11___mmap_ARPROT),
    .s01_axi_arqos(m_axi_rmem11___Stream2Mmap_11___mmap_ARQOS),
    .s01_axi_arready(m_axi_rmem11___Stream2Mmap_11___mmap_ARREADY),
    .s01_axi_arsize(m_axi_rmem11___Stream2Mmap_11___mmap_ARSIZE),
    .s01_axi_arvalid(m_axi_rmem11___Stream2Mmap_11___mmap_ARVALID),
    .s01_axi_awaddr(m_axi_rmem11___Stream2Mmap_11___mmap_AWADDR),
    .s01_axi_awburst(m_axi_rmem11___Stream2Mmap_11___mmap_AWBURST),
    .s01_axi_awcache(m_axi_rmem11___Stream2Mmap_11___mmap_AWCACHE),
    .s01_axi_awid(m_axi_rmem11___Stream2Mmap_11___mmap_AWID),
    .s01_axi_awlen(m_axi_rmem11___Stream2Mmap_11___mmap_AWLEN),
    .s01_axi_awlock(m_axi_rmem11___Stream2Mmap_11___mmap_AWLOCK),
    .s01_axi_awprot(m_axi_rmem11___Stream2Mmap_11___mmap_AWPROT),
    .s01_axi_awqos(m_axi_rmem11___Stream2Mmap_11___mmap_AWQOS),
    .s01_axi_awready(m_axi_rmem11___Stream2Mmap_11___mmap_AWREADY),
    .s01_axi_awsize(m_axi_rmem11___Stream2Mmap_11___mmap_AWSIZE),
    .s01_axi_awvalid(m_axi_rmem11___Stream2Mmap_11___mmap_AWVALID),
    .s01_axi_bid(m_axi_rmem11___Stream2Mmap_11___mmap_BID),
    .s01_axi_bready(m_axi_rmem11___Stream2Mmap_11___mmap_BREADY),
    .s01_axi_bresp(m_axi_rmem11___Stream2Mmap_11___mmap_BRESP),
    .s01_axi_bvalid(m_axi_rmem11___Stream2Mmap_11___mmap_BVALID),
    .s01_axi_rdata(m_axi_rmem11___Stream2Mmap_11___mmap_RDATA),
    .s01_axi_rid(m_axi_rmem11___Stream2Mmap_11___mmap_RID),
    .s01_axi_rlast(m_axi_rmem11___Stream2Mmap_11___mmap_RLAST),
    .s01_axi_rready(m_axi_rmem11___Stream2Mmap_11___mmap_RREADY),
    .s01_axi_rresp(m_axi_rmem11___Stream2Mmap_11___mmap_RRESP),
    .s01_axi_rvalid(m_axi_rmem11___Stream2Mmap_11___mmap_RVALID),
    .s01_axi_wdata(m_axi_rmem11___Stream2Mmap_11___mmap_WDATA),
    .s01_axi_wlast(m_axi_rmem11___Stream2Mmap_11___mmap_WLAST),
    .s01_axi_wready(m_axi_rmem11___Stream2Mmap_11___mmap_WREADY),
    .s01_axi_wstrb(m_axi_rmem11___Stream2Mmap_11___mmap_WSTRB),
    .s01_axi_wvalid(m_axi_rmem11___Stream2Mmap_11___mmap_WVALID)
  );


  (* keep_hierarchy = "yes" *) axi_crossbar_2x1
  #(
    .DATA_WIDTH(512),
    .ADDR_WIDTH(64),
    .S_ID_WIDTH(1),
    .M_ID_WIDTH(2),
    .M00_ADDR_WIDTH(64),
    .M00_ISSUE(16),
    .S00_THREADS(1),
    .S01_THREADS(1)
  )
  axi_crossbar_2x1__rmem12
  (
    .clk(ap_clk),
    .rst(ap_rst_n_inv),
    .m00_axi_araddr(m_axi_rmem12_ARADDR),
    .m00_axi_arburst(m_axi_rmem12_ARBURST),
    .m00_axi_arcache(m_axi_rmem12_ARCACHE),
    .m00_axi_arid(m_axi_rmem12_ARID),
    .m00_axi_arlen(m_axi_rmem12_ARLEN),
    .m00_axi_arlock(m_axi_rmem12_ARLOCK),
    .m00_axi_arprot(m_axi_rmem12_ARPROT),
    .m00_axi_arqos(m_axi_rmem12_ARQOS),
    .m00_axi_arready(m_axi_rmem12_ARREADY),
    .m00_axi_arsize(m_axi_rmem12_ARSIZE),
    .m00_axi_arvalid(m_axi_rmem12_ARVALID),
    .m00_axi_awaddr(m_axi_rmem12_AWADDR),
    .m00_axi_awburst(m_axi_rmem12_AWBURST),
    .m00_axi_awcache(m_axi_rmem12_AWCACHE),
    .m00_axi_awid(m_axi_rmem12_AWID),
    .m00_axi_awlen(m_axi_rmem12_AWLEN),
    .m00_axi_awlock(m_axi_rmem12_AWLOCK),
    .m00_axi_awprot(m_axi_rmem12_AWPROT),
    .m00_axi_awqos(m_axi_rmem12_AWQOS),
    .m00_axi_awready(m_axi_rmem12_AWREADY),
    .m00_axi_awsize(m_axi_rmem12_AWSIZE),
    .m00_axi_awvalid(m_axi_rmem12_AWVALID),
    .m00_axi_bid(m_axi_rmem12_BID),
    .m00_axi_bready(m_axi_rmem12_BREADY),
    .m00_axi_bresp(m_axi_rmem12_BRESP),
    .m00_axi_bvalid(m_axi_rmem12_BVALID),
    .m00_axi_rdata(m_axi_rmem12_RDATA),
    .m00_axi_rid(m_axi_rmem12_RID),
    .m00_axi_rlast(m_axi_rmem12_RLAST),
    .m00_axi_rready(m_axi_rmem12_RREADY),
    .m00_axi_rresp(m_axi_rmem12_RRESP),
    .m00_axi_rvalid(m_axi_rmem12_RVALID),
    .m00_axi_wdata(m_axi_rmem12_WDATA),
    .m00_axi_wlast(m_axi_rmem12_WLAST),
    .m00_axi_wready(m_axi_rmem12_WREADY),
    .m00_axi_wstrb(m_axi_rmem12_WSTRB),
    .m00_axi_wvalid(m_axi_rmem12_WVALID),
    .s00_axi_araddr(m_axi_rmem12___Mmap2Stream_12___mmap_ARADDR),
    .s00_axi_arburst(m_axi_rmem12___Mmap2Stream_12___mmap_ARBURST),
    .s00_axi_arcache(m_axi_rmem12___Mmap2Stream_12___mmap_ARCACHE),
    .s00_axi_arid(m_axi_rmem12___Mmap2Stream_12___mmap_ARID),
    .s00_axi_arlen(m_axi_rmem12___Mmap2Stream_12___mmap_ARLEN),
    .s00_axi_arlock(m_axi_rmem12___Mmap2Stream_12___mmap_ARLOCK),
    .s00_axi_arprot(m_axi_rmem12___Mmap2Stream_12___mmap_ARPROT),
    .s00_axi_arqos(m_axi_rmem12___Mmap2Stream_12___mmap_ARQOS),
    .s00_axi_arready(m_axi_rmem12___Mmap2Stream_12___mmap_ARREADY),
    .s00_axi_arsize(m_axi_rmem12___Mmap2Stream_12___mmap_ARSIZE),
    .s00_axi_arvalid(m_axi_rmem12___Mmap2Stream_12___mmap_ARVALID),
    .s00_axi_awaddr(m_axi_rmem12___Mmap2Stream_12___mmap_AWADDR),
    .s00_axi_awburst(m_axi_rmem12___Mmap2Stream_12___mmap_AWBURST),
    .s00_axi_awcache(m_axi_rmem12___Mmap2Stream_12___mmap_AWCACHE),
    .s00_axi_awid(m_axi_rmem12___Mmap2Stream_12___mmap_AWID),
    .s00_axi_awlen(m_axi_rmem12___Mmap2Stream_12___mmap_AWLEN),
    .s00_axi_awlock(m_axi_rmem12___Mmap2Stream_12___mmap_AWLOCK),
    .s00_axi_awprot(m_axi_rmem12___Mmap2Stream_12___mmap_AWPROT),
    .s00_axi_awqos(m_axi_rmem12___Mmap2Stream_12___mmap_AWQOS),
    .s00_axi_awready(m_axi_rmem12___Mmap2Stream_12___mmap_AWREADY),
    .s00_axi_awsize(m_axi_rmem12___Mmap2Stream_12___mmap_AWSIZE),
    .s00_axi_awvalid(m_axi_rmem12___Mmap2Stream_12___mmap_AWVALID),
    .s00_axi_bid(m_axi_rmem12___Mmap2Stream_12___mmap_BID),
    .s00_axi_bready(m_axi_rmem12___Mmap2Stream_12___mmap_BREADY),
    .s00_axi_bresp(m_axi_rmem12___Mmap2Stream_12___mmap_BRESP),
    .s00_axi_bvalid(m_axi_rmem12___Mmap2Stream_12___mmap_BVALID),
    .s00_axi_rdata(m_axi_rmem12___Mmap2Stream_12___mmap_RDATA),
    .s00_axi_rid(m_axi_rmem12___Mmap2Stream_12___mmap_RID),
    .s00_axi_rlast(m_axi_rmem12___Mmap2Stream_12___mmap_RLAST),
    .s00_axi_rready(m_axi_rmem12___Mmap2Stream_12___mmap_RREADY),
    .s00_axi_rresp(m_axi_rmem12___Mmap2Stream_12___mmap_RRESP),
    .s00_axi_rvalid(m_axi_rmem12___Mmap2Stream_12___mmap_RVALID),
    .s00_axi_wdata(m_axi_rmem12___Mmap2Stream_12___mmap_WDATA),
    .s00_axi_wlast(m_axi_rmem12___Mmap2Stream_12___mmap_WLAST),
    .s00_axi_wready(m_axi_rmem12___Mmap2Stream_12___mmap_WREADY),
    .s00_axi_wstrb(m_axi_rmem12___Mmap2Stream_12___mmap_WSTRB),
    .s00_axi_wvalid(m_axi_rmem12___Mmap2Stream_12___mmap_WVALID),
    .s01_axi_araddr(m_axi_rmem12___Stream2Mmap_12___mmap_ARADDR),
    .s01_axi_arburst(m_axi_rmem12___Stream2Mmap_12___mmap_ARBURST),
    .s01_axi_arcache(m_axi_rmem12___Stream2Mmap_12___mmap_ARCACHE),
    .s01_axi_arid(m_axi_rmem12___Stream2Mmap_12___mmap_ARID),
    .s01_axi_arlen(m_axi_rmem12___Stream2Mmap_12___mmap_ARLEN),
    .s01_axi_arlock(m_axi_rmem12___Stream2Mmap_12___mmap_ARLOCK),
    .s01_axi_arprot(m_axi_rmem12___Stream2Mmap_12___mmap_ARPROT),
    .s01_axi_arqos(m_axi_rmem12___Stream2Mmap_12___mmap_ARQOS),
    .s01_axi_arready(m_axi_rmem12___Stream2Mmap_12___mmap_ARREADY),
    .s01_axi_arsize(m_axi_rmem12___Stream2Mmap_12___mmap_ARSIZE),
    .s01_axi_arvalid(m_axi_rmem12___Stream2Mmap_12___mmap_ARVALID),
    .s01_axi_awaddr(m_axi_rmem12___Stream2Mmap_12___mmap_AWADDR),
    .s01_axi_awburst(m_axi_rmem12___Stream2Mmap_12___mmap_AWBURST),
    .s01_axi_awcache(m_axi_rmem12___Stream2Mmap_12___mmap_AWCACHE),
    .s01_axi_awid(m_axi_rmem12___Stream2Mmap_12___mmap_AWID),
    .s01_axi_awlen(m_axi_rmem12___Stream2Mmap_12___mmap_AWLEN),
    .s01_axi_awlock(m_axi_rmem12___Stream2Mmap_12___mmap_AWLOCK),
    .s01_axi_awprot(m_axi_rmem12___Stream2Mmap_12___mmap_AWPROT),
    .s01_axi_awqos(m_axi_rmem12___Stream2Mmap_12___mmap_AWQOS),
    .s01_axi_awready(m_axi_rmem12___Stream2Mmap_12___mmap_AWREADY),
    .s01_axi_awsize(m_axi_rmem12___Stream2Mmap_12___mmap_AWSIZE),
    .s01_axi_awvalid(m_axi_rmem12___Stream2Mmap_12___mmap_AWVALID),
    .s01_axi_bid(m_axi_rmem12___Stream2Mmap_12___mmap_BID),
    .s01_axi_bready(m_axi_rmem12___Stream2Mmap_12___mmap_BREADY),
    .s01_axi_bresp(m_axi_rmem12___Stream2Mmap_12___mmap_BRESP),
    .s01_axi_bvalid(m_axi_rmem12___Stream2Mmap_12___mmap_BVALID),
    .s01_axi_rdata(m_axi_rmem12___Stream2Mmap_12___mmap_RDATA),
    .s01_axi_rid(m_axi_rmem12___Stream2Mmap_12___mmap_RID),
    .s01_axi_rlast(m_axi_rmem12___Stream2Mmap_12___mmap_RLAST),
    .s01_axi_rready(m_axi_rmem12___Stream2Mmap_12___mmap_RREADY),
    .s01_axi_rresp(m_axi_rmem12___Stream2Mmap_12___mmap_RRESP),
    .s01_axi_rvalid(m_axi_rmem12___Stream2Mmap_12___mmap_RVALID),
    .s01_axi_wdata(m_axi_rmem12___Stream2Mmap_12___mmap_WDATA),
    .s01_axi_wlast(m_axi_rmem12___Stream2Mmap_12___mmap_WLAST),
    .s01_axi_wready(m_axi_rmem12___Stream2Mmap_12___mmap_WREADY),
    .s01_axi_wstrb(m_axi_rmem12___Stream2Mmap_12___mmap_WSTRB),
    .s01_axi_wvalid(m_axi_rmem12___Stream2Mmap_12___mmap_WVALID)
  );


  (* keep_hierarchy = "yes" *) axi_crossbar_2x1
  #(
    .DATA_WIDTH(512),
    .ADDR_WIDTH(64),
    .S_ID_WIDTH(1),
    .M_ID_WIDTH(2),
    .M00_ADDR_WIDTH(64),
    .M00_ISSUE(16),
    .S00_THREADS(1),
    .S01_THREADS(1)
  )
  axi_crossbar_2x1__rmem13
  (
    .clk(ap_clk),
    .rst(ap_rst_n_inv),
    .m00_axi_araddr(m_axi_rmem13_ARADDR),
    .m00_axi_arburst(m_axi_rmem13_ARBURST),
    .m00_axi_arcache(m_axi_rmem13_ARCACHE),
    .m00_axi_arid(m_axi_rmem13_ARID),
    .m00_axi_arlen(m_axi_rmem13_ARLEN),
    .m00_axi_arlock(m_axi_rmem13_ARLOCK),
    .m00_axi_arprot(m_axi_rmem13_ARPROT),
    .m00_axi_arqos(m_axi_rmem13_ARQOS),
    .m00_axi_arready(m_axi_rmem13_ARREADY),
    .m00_axi_arsize(m_axi_rmem13_ARSIZE),
    .m00_axi_arvalid(m_axi_rmem13_ARVALID),
    .m00_axi_awaddr(m_axi_rmem13_AWADDR),
    .m00_axi_awburst(m_axi_rmem13_AWBURST),
    .m00_axi_awcache(m_axi_rmem13_AWCACHE),
    .m00_axi_awid(m_axi_rmem13_AWID),
    .m00_axi_awlen(m_axi_rmem13_AWLEN),
    .m00_axi_awlock(m_axi_rmem13_AWLOCK),
    .m00_axi_awprot(m_axi_rmem13_AWPROT),
    .m00_axi_awqos(m_axi_rmem13_AWQOS),
    .m00_axi_awready(m_axi_rmem13_AWREADY),
    .m00_axi_awsize(m_axi_rmem13_AWSIZE),
    .m00_axi_awvalid(m_axi_rmem13_AWVALID),
    .m00_axi_bid(m_axi_rmem13_BID),
    .m00_axi_bready(m_axi_rmem13_BREADY),
    .m00_axi_bresp(m_axi_rmem13_BRESP),
    .m00_axi_bvalid(m_axi_rmem13_BVALID),
    .m00_axi_rdata(m_axi_rmem13_RDATA),
    .m00_axi_rid(m_axi_rmem13_RID),
    .m00_axi_rlast(m_axi_rmem13_RLAST),
    .m00_axi_rready(m_axi_rmem13_RREADY),
    .m00_axi_rresp(m_axi_rmem13_RRESP),
    .m00_axi_rvalid(m_axi_rmem13_RVALID),
    .m00_axi_wdata(m_axi_rmem13_WDATA),
    .m00_axi_wlast(m_axi_rmem13_WLAST),
    .m00_axi_wready(m_axi_rmem13_WREADY),
    .m00_axi_wstrb(m_axi_rmem13_WSTRB),
    .m00_axi_wvalid(m_axi_rmem13_WVALID),
    .s00_axi_araddr(m_axi_rmem13___Mmap2Stream_13___mmap_ARADDR),
    .s00_axi_arburst(m_axi_rmem13___Mmap2Stream_13___mmap_ARBURST),
    .s00_axi_arcache(m_axi_rmem13___Mmap2Stream_13___mmap_ARCACHE),
    .s00_axi_arid(m_axi_rmem13___Mmap2Stream_13___mmap_ARID),
    .s00_axi_arlen(m_axi_rmem13___Mmap2Stream_13___mmap_ARLEN),
    .s00_axi_arlock(m_axi_rmem13___Mmap2Stream_13___mmap_ARLOCK),
    .s00_axi_arprot(m_axi_rmem13___Mmap2Stream_13___mmap_ARPROT),
    .s00_axi_arqos(m_axi_rmem13___Mmap2Stream_13___mmap_ARQOS),
    .s00_axi_arready(m_axi_rmem13___Mmap2Stream_13___mmap_ARREADY),
    .s00_axi_arsize(m_axi_rmem13___Mmap2Stream_13___mmap_ARSIZE),
    .s00_axi_arvalid(m_axi_rmem13___Mmap2Stream_13___mmap_ARVALID),
    .s00_axi_awaddr(m_axi_rmem13___Mmap2Stream_13___mmap_AWADDR),
    .s00_axi_awburst(m_axi_rmem13___Mmap2Stream_13___mmap_AWBURST),
    .s00_axi_awcache(m_axi_rmem13___Mmap2Stream_13___mmap_AWCACHE),
    .s00_axi_awid(m_axi_rmem13___Mmap2Stream_13___mmap_AWID),
    .s00_axi_awlen(m_axi_rmem13___Mmap2Stream_13___mmap_AWLEN),
    .s00_axi_awlock(m_axi_rmem13___Mmap2Stream_13___mmap_AWLOCK),
    .s00_axi_awprot(m_axi_rmem13___Mmap2Stream_13___mmap_AWPROT),
    .s00_axi_awqos(m_axi_rmem13___Mmap2Stream_13___mmap_AWQOS),
    .s00_axi_awready(m_axi_rmem13___Mmap2Stream_13___mmap_AWREADY),
    .s00_axi_awsize(m_axi_rmem13___Mmap2Stream_13___mmap_AWSIZE),
    .s00_axi_awvalid(m_axi_rmem13___Mmap2Stream_13___mmap_AWVALID),
    .s00_axi_bid(m_axi_rmem13___Mmap2Stream_13___mmap_BID),
    .s00_axi_bready(m_axi_rmem13___Mmap2Stream_13___mmap_BREADY),
    .s00_axi_bresp(m_axi_rmem13___Mmap2Stream_13___mmap_BRESP),
    .s00_axi_bvalid(m_axi_rmem13___Mmap2Stream_13___mmap_BVALID),
    .s00_axi_rdata(m_axi_rmem13___Mmap2Stream_13___mmap_RDATA),
    .s00_axi_rid(m_axi_rmem13___Mmap2Stream_13___mmap_RID),
    .s00_axi_rlast(m_axi_rmem13___Mmap2Stream_13___mmap_RLAST),
    .s00_axi_rready(m_axi_rmem13___Mmap2Stream_13___mmap_RREADY),
    .s00_axi_rresp(m_axi_rmem13___Mmap2Stream_13___mmap_RRESP),
    .s00_axi_rvalid(m_axi_rmem13___Mmap2Stream_13___mmap_RVALID),
    .s00_axi_wdata(m_axi_rmem13___Mmap2Stream_13___mmap_WDATA),
    .s00_axi_wlast(m_axi_rmem13___Mmap2Stream_13___mmap_WLAST),
    .s00_axi_wready(m_axi_rmem13___Mmap2Stream_13___mmap_WREADY),
    .s00_axi_wstrb(m_axi_rmem13___Mmap2Stream_13___mmap_WSTRB),
    .s00_axi_wvalid(m_axi_rmem13___Mmap2Stream_13___mmap_WVALID),
    .s01_axi_araddr(m_axi_rmem13___Stream2Mmap_13___mmap_ARADDR),
    .s01_axi_arburst(m_axi_rmem13___Stream2Mmap_13___mmap_ARBURST),
    .s01_axi_arcache(m_axi_rmem13___Stream2Mmap_13___mmap_ARCACHE),
    .s01_axi_arid(m_axi_rmem13___Stream2Mmap_13___mmap_ARID),
    .s01_axi_arlen(m_axi_rmem13___Stream2Mmap_13___mmap_ARLEN),
    .s01_axi_arlock(m_axi_rmem13___Stream2Mmap_13___mmap_ARLOCK),
    .s01_axi_arprot(m_axi_rmem13___Stream2Mmap_13___mmap_ARPROT),
    .s01_axi_arqos(m_axi_rmem13___Stream2Mmap_13___mmap_ARQOS),
    .s01_axi_arready(m_axi_rmem13___Stream2Mmap_13___mmap_ARREADY),
    .s01_axi_arsize(m_axi_rmem13___Stream2Mmap_13___mmap_ARSIZE),
    .s01_axi_arvalid(m_axi_rmem13___Stream2Mmap_13___mmap_ARVALID),
    .s01_axi_awaddr(m_axi_rmem13___Stream2Mmap_13___mmap_AWADDR),
    .s01_axi_awburst(m_axi_rmem13___Stream2Mmap_13___mmap_AWBURST),
    .s01_axi_awcache(m_axi_rmem13___Stream2Mmap_13___mmap_AWCACHE),
    .s01_axi_awid(m_axi_rmem13___Stream2Mmap_13___mmap_AWID),
    .s01_axi_awlen(m_axi_rmem13___Stream2Mmap_13___mmap_AWLEN),
    .s01_axi_awlock(m_axi_rmem13___Stream2Mmap_13___mmap_AWLOCK),
    .s01_axi_awprot(m_axi_rmem13___Stream2Mmap_13___mmap_AWPROT),
    .s01_axi_awqos(m_axi_rmem13___Stream2Mmap_13___mmap_AWQOS),
    .s01_axi_awready(m_axi_rmem13___Stream2Mmap_13___mmap_AWREADY),
    .s01_axi_awsize(m_axi_rmem13___Stream2Mmap_13___mmap_AWSIZE),
    .s01_axi_awvalid(m_axi_rmem13___Stream2Mmap_13___mmap_AWVALID),
    .s01_axi_bid(m_axi_rmem13___Stream2Mmap_13___mmap_BID),
    .s01_axi_bready(m_axi_rmem13___Stream2Mmap_13___mmap_BREADY),
    .s01_axi_bresp(m_axi_rmem13___Stream2Mmap_13___mmap_BRESP),
    .s01_axi_bvalid(m_axi_rmem13___Stream2Mmap_13___mmap_BVALID),
    .s01_axi_rdata(m_axi_rmem13___Stream2Mmap_13___mmap_RDATA),
    .s01_axi_rid(m_axi_rmem13___Stream2Mmap_13___mmap_RID),
    .s01_axi_rlast(m_axi_rmem13___Stream2Mmap_13___mmap_RLAST),
    .s01_axi_rready(m_axi_rmem13___Stream2Mmap_13___mmap_RREADY),
    .s01_axi_rresp(m_axi_rmem13___Stream2Mmap_13___mmap_RRESP),
    .s01_axi_rvalid(m_axi_rmem13___Stream2Mmap_13___mmap_RVALID),
    .s01_axi_wdata(m_axi_rmem13___Stream2Mmap_13___mmap_WDATA),
    .s01_axi_wlast(m_axi_rmem13___Stream2Mmap_13___mmap_WLAST),
    .s01_axi_wready(m_axi_rmem13___Stream2Mmap_13___mmap_WREADY),
    .s01_axi_wstrb(m_axi_rmem13___Stream2Mmap_13___mmap_WSTRB),
    .s01_axi_wvalid(m_axi_rmem13___Stream2Mmap_13___mmap_WVALID)
  );


  (* keep_hierarchy = "yes" *) axi_crossbar_2x1
  #(
    .DATA_WIDTH(512),
    .ADDR_WIDTH(64),
    .S_ID_WIDTH(1),
    .M_ID_WIDTH(2),
    .M00_ADDR_WIDTH(64),
    .M00_ISSUE(16),
    .S00_THREADS(1),
    .S01_THREADS(1)
  )
  axi_crossbar_2x1__rmem14
  (
    .clk(ap_clk),
    .rst(ap_rst_n_inv),
    .m00_axi_araddr(m_axi_rmem14_ARADDR),
    .m00_axi_arburst(m_axi_rmem14_ARBURST),
    .m00_axi_arcache(m_axi_rmem14_ARCACHE),
    .m00_axi_arid(m_axi_rmem14_ARID),
    .m00_axi_arlen(m_axi_rmem14_ARLEN),
    .m00_axi_arlock(m_axi_rmem14_ARLOCK),
    .m00_axi_arprot(m_axi_rmem14_ARPROT),
    .m00_axi_arqos(m_axi_rmem14_ARQOS),
    .m00_axi_arready(m_axi_rmem14_ARREADY),
    .m00_axi_arsize(m_axi_rmem14_ARSIZE),
    .m00_axi_arvalid(m_axi_rmem14_ARVALID),
    .m00_axi_awaddr(m_axi_rmem14_AWADDR),
    .m00_axi_awburst(m_axi_rmem14_AWBURST),
    .m00_axi_awcache(m_axi_rmem14_AWCACHE),
    .m00_axi_awid(m_axi_rmem14_AWID),
    .m00_axi_awlen(m_axi_rmem14_AWLEN),
    .m00_axi_awlock(m_axi_rmem14_AWLOCK),
    .m00_axi_awprot(m_axi_rmem14_AWPROT),
    .m00_axi_awqos(m_axi_rmem14_AWQOS),
    .m00_axi_awready(m_axi_rmem14_AWREADY),
    .m00_axi_awsize(m_axi_rmem14_AWSIZE),
    .m00_axi_awvalid(m_axi_rmem14_AWVALID),
    .m00_axi_bid(m_axi_rmem14_BID),
    .m00_axi_bready(m_axi_rmem14_BREADY),
    .m00_axi_bresp(m_axi_rmem14_BRESP),
    .m00_axi_bvalid(m_axi_rmem14_BVALID),
    .m00_axi_rdata(m_axi_rmem14_RDATA),
    .m00_axi_rid(m_axi_rmem14_RID),
    .m00_axi_rlast(m_axi_rmem14_RLAST),
    .m00_axi_rready(m_axi_rmem14_RREADY),
    .m00_axi_rresp(m_axi_rmem14_RRESP),
    .m00_axi_rvalid(m_axi_rmem14_RVALID),
    .m00_axi_wdata(m_axi_rmem14_WDATA),
    .m00_axi_wlast(m_axi_rmem14_WLAST),
    .m00_axi_wready(m_axi_rmem14_WREADY),
    .m00_axi_wstrb(m_axi_rmem14_WSTRB),
    .m00_axi_wvalid(m_axi_rmem14_WVALID),
    .s00_axi_araddr(m_axi_rmem14___Mmap2Stream_14___mmap_ARADDR),
    .s00_axi_arburst(m_axi_rmem14___Mmap2Stream_14___mmap_ARBURST),
    .s00_axi_arcache(m_axi_rmem14___Mmap2Stream_14___mmap_ARCACHE),
    .s00_axi_arid(m_axi_rmem14___Mmap2Stream_14___mmap_ARID),
    .s00_axi_arlen(m_axi_rmem14___Mmap2Stream_14___mmap_ARLEN),
    .s00_axi_arlock(m_axi_rmem14___Mmap2Stream_14___mmap_ARLOCK),
    .s00_axi_arprot(m_axi_rmem14___Mmap2Stream_14___mmap_ARPROT),
    .s00_axi_arqos(m_axi_rmem14___Mmap2Stream_14___mmap_ARQOS),
    .s00_axi_arready(m_axi_rmem14___Mmap2Stream_14___mmap_ARREADY),
    .s00_axi_arsize(m_axi_rmem14___Mmap2Stream_14___mmap_ARSIZE),
    .s00_axi_arvalid(m_axi_rmem14___Mmap2Stream_14___mmap_ARVALID),
    .s00_axi_awaddr(m_axi_rmem14___Mmap2Stream_14___mmap_AWADDR),
    .s00_axi_awburst(m_axi_rmem14___Mmap2Stream_14___mmap_AWBURST),
    .s00_axi_awcache(m_axi_rmem14___Mmap2Stream_14___mmap_AWCACHE),
    .s00_axi_awid(m_axi_rmem14___Mmap2Stream_14___mmap_AWID),
    .s00_axi_awlen(m_axi_rmem14___Mmap2Stream_14___mmap_AWLEN),
    .s00_axi_awlock(m_axi_rmem14___Mmap2Stream_14___mmap_AWLOCK),
    .s00_axi_awprot(m_axi_rmem14___Mmap2Stream_14___mmap_AWPROT),
    .s00_axi_awqos(m_axi_rmem14___Mmap2Stream_14___mmap_AWQOS),
    .s00_axi_awready(m_axi_rmem14___Mmap2Stream_14___mmap_AWREADY),
    .s00_axi_awsize(m_axi_rmem14___Mmap2Stream_14___mmap_AWSIZE),
    .s00_axi_awvalid(m_axi_rmem14___Mmap2Stream_14___mmap_AWVALID),
    .s00_axi_bid(m_axi_rmem14___Mmap2Stream_14___mmap_BID),
    .s00_axi_bready(m_axi_rmem14___Mmap2Stream_14___mmap_BREADY),
    .s00_axi_bresp(m_axi_rmem14___Mmap2Stream_14___mmap_BRESP),
    .s00_axi_bvalid(m_axi_rmem14___Mmap2Stream_14___mmap_BVALID),
    .s00_axi_rdata(m_axi_rmem14___Mmap2Stream_14___mmap_RDATA),
    .s00_axi_rid(m_axi_rmem14___Mmap2Stream_14___mmap_RID),
    .s00_axi_rlast(m_axi_rmem14___Mmap2Stream_14___mmap_RLAST),
    .s00_axi_rready(m_axi_rmem14___Mmap2Stream_14___mmap_RREADY),
    .s00_axi_rresp(m_axi_rmem14___Mmap2Stream_14___mmap_RRESP),
    .s00_axi_rvalid(m_axi_rmem14___Mmap2Stream_14___mmap_RVALID),
    .s00_axi_wdata(m_axi_rmem14___Mmap2Stream_14___mmap_WDATA),
    .s00_axi_wlast(m_axi_rmem14___Mmap2Stream_14___mmap_WLAST),
    .s00_axi_wready(m_axi_rmem14___Mmap2Stream_14___mmap_WREADY),
    .s00_axi_wstrb(m_axi_rmem14___Mmap2Stream_14___mmap_WSTRB),
    .s00_axi_wvalid(m_axi_rmem14___Mmap2Stream_14___mmap_WVALID),
    .s01_axi_araddr(m_axi_rmem14___Stream2Mmap_14___mmap_ARADDR),
    .s01_axi_arburst(m_axi_rmem14___Stream2Mmap_14___mmap_ARBURST),
    .s01_axi_arcache(m_axi_rmem14___Stream2Mmap_14___mmap_ARCACHE),
    .s01_axi_arid(m_axi_rmem14___Stream2Mmap_14___mmap_ARID),
    .s01_axi_arlen(m_axi_rmem14___Stream2Mmap_14___mmap_ARLEN),
    .s01_axi_arlock(m_axi_rmem14___Stream2Mmap_14___mmap_ARLOCK),
    .s01_axi_arprot(m_axi_rmem14___Stream2Mmap_14___mmap_ARPROT),
    .s01_axi_arqos(m_axi_rmem14___Stream2Mmap_14___mmap_ARQOS),
    .s01_axi_arready(m_axi_rmem14___Stream2Mmap_14___mmap_ARREADY),
    .s01_axi_arsize(m_axi_rmem14___Stream2Mmap_14___mmap_ARSIZE),
    .s01_axi_arvalid(m_axi_rmem14___Stream2Mmap_14___mmap_ARVALID),
    .s01_axi_awaddr(m_axi_rmem14___Stream2Mmap_14___mmap_AWADDR),
    .s01_axi_awburst(m_axi_rmem14___Stream2Mmap_14___mmap_AWBURST),
    .s01_axi_awcache(m_axi_rmem14___Stream2Mmap_14___mmap_AWCACHE),
    .s01_axi_awid(m_axi_rmem14___Stream2Mmap_14___mmap_AWID),
    .s01_axi_awlen(m_axi_rmem14___Stream2Mmap_14___mmap_AWLEN),
    .s01_axi_awlock(m_axi_rmem14___Stream2Mmap_14___mmap_AWLOCK),
    .s01_axi_awprot(m_axi_rmem14___Stream2Mmap_14___mmap_AWPROT),
    .s01_axi_awqos(m_axi_rmem14___Stream2Mmap_14___mmap_AWQOS),
    .s01_axi_awready(m_axi_rmem14___Stream2Mmap_14___mmap_AWREADY),
    .s01_axi_awsize(m_axi_rmem14___Stream2Mmap_14___mmap_AWSIZE),
    .s01_axi_awvalid(m_axi_rmem14___Stream2Mmap_14___mmap_AWVALID),
    .s01_axi_bid(m_axi_rmem14___Stream2Mmap_14___mmap_BID),
    .s01_axi_bready(m_axi_rmem14___Stream2Mmap_14___mmap_BREADY),
    .s01_axi_bresp(m_axi_rmem14___Stream2Mmap_14___mmap_BRESP),
    .s01_axi_bvalid(m_axi_rmem14___Stream2Mmap_14___mmap_BVALID),
    .s01_axi_rdata(m_axi_rmem14___Stream2Mmap_14___mmap_RDATA),
    .s01_axi_rid(m_axi_rmem14___Stream2Mmap_14___mmap_RID),
    .s01_axi_rlast(m_axi_rmem14___Stream2Mmap_14___mmap_RLAST),
    .s01_axi_rready(m_axi_rmem14___Stream2Mmap_14___mmap_RREADY),
    .s01_axi_rresp(m_axi_rmem14___Stream2Mmap_14___mmap_RRESP),
    .s01_axi_rvalid(m_axi_rmem14___Stream2Mmap_14___mmap_RVALID),
    .s01_axi_wdata(m_axi_rmem14___Stream2Mmap_14___mmap_WDATA),
    .s01_axi_wlast(m_axi_rmem14___Stream2Mmap_14___mmap_WLAST),
    .s01_axi_wready(m_axi_rmem14___Stream2Mmap_14___mmap_WREADY),
    .s01_axi_wstrb(m_axi_rmem14___Stream2Mmap_14___mmap_WSTRB),
    .s01_axi_wvalid(m_axi_rmem14___Stream2Mmap_14___mmap_WVALID)
  );


  (* keep_hierarchy = "yes" *) axi_crossbar_2x1
  #(
    .DATA_WIDTH(512),
    .ADDR_WIDTH(64),
    .S_ID_WIDTH(1),
    .M_ID_WIDTH(2),
    .M00_ADDR_WIDTH(64),
    .M00_ISSUE(16),
    .S00_THREADS(1),
    .S01_THREADS(1)
  )
  axi_crossbar_2x1__rmem15
  (
    .clk(ap_clk),
    .rst(ap_rst_n_inv),
    .m00_axi_araddr(m_axi_rmem15_ARADDR),
    .m00_axi_arburst(m_axi_rmem15_ARBURST),
    .m00_axi_arcache(m_axi_rmem15_ARCACHE),
    .m00_axi_arid(m_axi_rmem15_ARID),
    .m00_axi_arlen(m_axi_rmem15_ARLEN),
    .m00_axi_arlock(m_axi_rmem15_ARLOCK),
    .m00_axi_arprot(m_axi_rmem15_ARPROT),
    .m00_axi_arqos(m_axi_rmem15_ARQOS),
    .m00_axi_arready(m_axi_rmem15_ARREADY),
    .m00_axi_arsize(m_axi_rmem15_ARSIZE),
    .m00_axi_arvalid(m_axi_rmem15_ARVALID),
    .m00_axi_awaddr(m_axi_rmem15_AWADDR),
    .m00_axi_awburst(m_axi_rmem15_AWBURST),
    .m00_axi_awcache(m_axi_rmem15_AWCACHE),
    .m00_axi_awid(m_axi_rmem15_AWID),
    .m00_axi_awlen(m_axi_rmem15_AWLEN),
    .m00_axi_awlock(m_axi_rmem15_AWLOCK),
    .m00_axi_awprot(m_axi_rmem15_AWPROT),
    .m00_axi_awqos(m_axi_rmem15_AWQOS),
    .m00_axi_awready(m_axi_rmem15_AWREADY),
    .m00_axi_awsize(m_axi_rmem15_AWSIZE),
    .m00_axi_awvalid(m_axi_rmem15_AWVALID),
    .m00_axi_bid(m_axi_rmem15_BID),
    .m00_axi_bready(m_axi_rmem15_BREADY),
    .m00_axi_bresp(m_axi_rmem15_BRESP),
    .m00_axi_bvalid(m_axi_rmem15_BVALID),
    .m00_axi_rdata(m_axi_rmem15_RDATA),
    .m00_axi_rid(m_axi_rmem15_RID),
    .m00_axi_rlast(m_axi_rmem15_RLAST),
    .m00_axi_rready(m_axi_rmem15_RREADY),
    .m00_axi_rresp(m_axi_rmem15_RRESP),
    .m00_axi_rvalid(m_axi_rmem15_RVALID),
    .m00_axi_wdata(m_axi_rmem15_WDATA),
    .m00_axi_wlast(m_axi_rmem15_WLAST),
    .m00_axi_wready(m_axi_rmem15_WREADY),
    .m00_axi_wstrb(m_axi_rmem15_WSTRB),
    .m00_axi_wvalid(m_axi_rmem15_WVALID),
    .s00_axi_araddr(m_axi_rmem15___Mmap2Stream_15___mmap_ARADDR),
    .s00_axi_arburst(m_axi_rmem15___Mmap2Stream_15___mmap_ARBURST),
    .s00_axi_arcache(m_axi_rmem15___Mmap2Stream_15___mmap_ARCACHE),
    .s00_axi_arid(m_axi_rmem15___Mmap2Stream_15___mmap_ARID),
    .s00_axi_arlen(m_axi_rmem15___Mmap2Stream_15___mmap_ARLEN),
    .s00_axi_arlock(m_axi_rmem15___Mmap2Stream_15___mmap_ARLOCK),
    .s00_axi_arprot(m_axi_rmem15___Mmap2Stream_15___mmap_ARPROT),
    .s00_axi_arqos(m_axi_rmem15___Mmap2Stream_15___mmap_ARQOS),
    .s00_axi_arready(m_axi_rmem15___Mmap2Stream_15___mmap_ARREADY),
    .s00_axi_arsize(m_axi_rmem15___Mmap2Stream_15___mmap_ARSIZE),
    .s00_axi_arvalid(m_axi_rmem15___Mmap2Stream_15___mmap_ARVALID),
    .s00_axi_awaddr(m_axi_rmem15___Mmap2Stream_15___mmap_AWADDR),
    .s00_axi_awburst(m_axi_rmem15___Mmap2Stream_15___mmap_AWBURST),
    .s00_axi_awcache(m_axi_rmem15___Mmap2Stream_15___mmap_AWCACHE),
    .s00_axi_awid(m_axi_rmem15___Mmap2Stream_15___mmap_AWID),
    .s00_axi_awlen(m_axi_rmem15___Mmap2Stream_15___mmap_AWLEN),
    .s00_axi_awlock(m_axi_rmem15___Mmap2Stream_15___mmap_AWLOCK),
    .s00_axi_awprot(m_axi_rmem15___Mmap2Stream_15___mmap_AWPROT),
    .s00_axi_awqos(m_axi_rmem15___Mmap2Stream_15___mmap_AWQOS),
    .s00_axi_awready(m_axi_rmem15___Mmap2Stream_15___mmap_AWREADY),
    .s00_axi_awsize(m_axi_rmem15___Mmap2Stream_15___mmap_AWSIZE),
    .s00_axi_awvalid(m_axi_rmem15___Mmap2Stream_15___mmap_AWVALID),
    .s00_axi_bid(m_axi_rmem15___Mmap2Stream_15___mmap_BID),
    .s00_axi_bready(m_axi_rmem15___Mmap2Stream_15___mmap_BREADY),
    .s00_axi_bresp(m_axi_rmem15___Mmap2Stream_15___mmap_BRESP),
    .s00_axi_bvalid(m_axi_rmem15___Mmap2Stream_15___mmap_BVALID),
    .s00_axi_rdata(m_axi_rmem15___Mmap2Stream_15___mmap_RDATA),
    .s00_axi_rid(m_axi_rmem15___Mmap2Stream_15___mmap_RID),
    .s00_axi_rlast(m_axi_rmem15___Mmap2Stream_15___mmap_RLAST),
    .s00_axi_rready(m_axi_rmem15___Mmap2Stream_15___mmap_RREADY),
    .s00_axi_rresp(m_axi_rmem15___Mmap2Stream_15___mmap_RRESP),
    .s00_axi_rvalid(m_axi_rmem15___Mmap2Stream_15___mmap_RVALID),
    .s00_axi_wdata(m_axi_rmem15___Mmap2Stream_15___mmap_WDATA),
    .s00_axi_wlast(m_axi_rmem15___Mmap2Stream_15___mmap_WLAST),
    .s00_axi_wready(m_axi_rmem15___Mmap2Stream_15___mmap_WREADY),
    .s00_axi_wstrb(m_axi_rmem15___Mmap2Stream_15___mmap_WSTRB),
    .s00_axi_wvalid(m_axi_rmem15___Mmap2Stream_15___mmap_WVALID),
    .s01_axi_araddr(m_axi_rmem15___Stream2Mmap_15___mmap_ARADDR),
    .s01_axi_arburst(m_axi_rmem15___Stream2Mmap_15___mmap_ARBURST),
    .s01_axi_arcache(m_axi_rmem15___Stream2Mmap_15___mmap_ARCACHE),
    .s01_axi_arid(m_axi_rmem15___Stream2Mmap_15___mmap_ARID),
    .s01_axi_arlen(m_axi_rmem15___Stream2Mmap_15___mmap_ARLEN),
    .s01_axi_arlock(m_axi_rmem15___Stream2Mmap_15___mmap_ARLOCK),
    .s01_axi_arprot(m_axi_rmem15___Stream2Mmap_15___mmap_ARPROT),
    .s01_axi_arqos(m_axi_rmem15___Stream2Mmap_15___mmap_ARQOS),
    .s01_axi_arready(m_axi_rmem15___Stream2Mmap_15___mmap_ARREADY),
    .s01_axi_arsize(m_axi_rmem15___Stream2Mmap_15___mmap_ARSIZE),
    .s01_axi_arvalid(m_axi_rmem15___Stream2Mmap_15___mmap_ARVALID),
    .s01_axi_awaddr(m_axi_rmem15___Stream2Mmap_15___mmap_AWADDR),
    .s01_axi_awburst(m_axi_rmem15___Stream2Mmap_15___mmap_AWBURST),
    .s01_axi_awcache(m_axi_rmem15___Stream2Mmap_15___mmap_AWCACHE),
    .s01_axi_awid(m_axi_rmem15___Stream2Mmap_15___mmap_AWID),
    .s01_axi_awlen(m_axi_rmem15___Stream2Mmap_15___mmap_AWLEN),
    .s01_axi_awlock(m_axi_rmem15___Stream2Mmap_15___mmap_AWLOCK),
    .s01_axi_awprot(m_axi_rmem15___Stream2Mmap_15___mmap_AWPROT),
    .s01_axi_awqos(m_axi_rmem15___Stream2Mmap_15___mmap_AWQOS),
    .s01_axi_awready(m_axi_rmem15___Stream2Mmap_15___mmap_AWREADY),
    .s01_axi_awsize(m_axi_rmem15___Stream2Mmap_15___mmap_AWSIZE),
    .s01_axi_awvalid(m_axi_rmem15___Stream2Mmap_15___mmap_AWVALID),
    .s01_axi_bid(m_axi_rmem15___Stream2Mmap_15___mmap_BID),
    .s01_axi_bready(m_axi_rmem15___Stream2Mmap_15___mmap_BREADY),
    .s01_axi_bresp(m_axi_rmem15___Stream2Mmap_15___mmap_BRESP),
    .s01_axi_bvalid(m_axi_rmem15___Stream2Mmap_15___mmap_BVALID),
    .s01_axi_rdata(m_axi_rmem15___Stream2Mmap_15___mmap_RDATA),
    .s01_axi_rid(m_axi_rmem15___Stream2Mmap_15___mmap_RID),
    .s01_axi_rlast(m_axi_rmem15___Stream2Mmap_15___mmap_RLAST),
    .s01_axi_rready(m_axi_rmem15___Stream2Mmap_15___mmap_RREADY),
    .s01_axi_rresp(m_axi_rmem15___Stream2Mmap_15___mmap_RRESP),
    .s01_axi_rvalid(m_axi_rmem15___Stream2Mmap_15___mmap_RVALID),
    .s01_axi_wdata(m_axi_rmem15___Stream2Mmap_15___mmap_WDATA),
    .s01_axi_wlast(m_axi_rmem15___Stream2Mmap_15___mmap_WLAST),
    .s01_axi_wready(m_axi_rmem15___Stream2Mmap_15___mmap_WREADY),
    .s01_axi_wstrb(m_axi_rmem15___Stream2Mmap_15___mmap_WSTRB),
    .s01_axi_wvalid(m_axi_rmem15___Stream2Mmap_15___mmap_WVALID)
  );


  (* keep_hierarchy = "yes" *) axi_crossbar_2x1
  #(
    .DATA_WIDTH(512),
    .ADDR_WIDTH(64),
    .S_ID_WIDTH(1),
    .M_ID_WIDTH(2),
    .M00_ADDR_WIDTH(64),
    .M00_ISSUE(16),
    .S00_THREADS(1),
    .S01_THREADS(1)
  )
  axi_crossbar_2x1__rmem16
  (
    .clk(ap_clk),
    .rst(ap_rst_n_inv),
    .m00_axi_araddr(m_axi_rmem16_ARADDR),
    .m00_axi_arburst(m_axi_rmem16_ARBURST),
    .m00_axi_arcache(m_axi_rmem16_ARCACHE),
    .m00_axi_arid(m_axi_rmem16_ARID),
    .m00_axi_arlen(m_axi_rmem16_ARLEN),
    .m00_axi_arlock(m_axi_rmem16_ARLOCK),
    .m00_axi_arprot(m_axi_rmem16_ARPROT),
    .m00_axi_arqos(m_axi_rmem16_ARQOS),
    .m00_axi_arready(m_axi_rmem16_ARREADY),
    .m00_axi_arsize(m_axi_rmem16_ARSIZE),
    .m00_axi_arvalid(m_axi_rmem16_ARVALID),
    .m00_axi_awaddr(m_axi_rmem16_AWADDR),
    .m00_axi_awburst(m_axi_rmem16_AWBURST),
    .m00_axi_awcache(m_axi_rmem16_AWCACHE),
    .m00_axi_awid(m_axi_rmem16_AWID),
    .m00_axi_awlen(m_axi_rmem16_AWLEN),
    .m00_axi_awlock(m_axi_rmem16_AWLOCK),
    .m00_axi_awprot(m_axi_rmem16_AWPROT),
    .m00_axi_awqos(m_axi_rmem16_AWQOS),
    .m00_axi_awready(m_axi_rmem16_AWREADY),
    .m00_axi_awsize(m_axi_rmem16_AWSIZE),
    .m00_axi_awvalid(m_axi_rmem16_AWVALID),
    .m00_axi_bid(m_axi_rmem16_BID),
    .m00_axi_bready(m_axi_rmem16_BREADY),
    .m00_axi_bresp(m_axi_rmem16_BRESP),
    .m00_axi_bvalid(m_axi_rmem16_BVALID),
    .m00_axi_rdata(m_axi_rmem16_RDATA),
    .m00_axi_rid(m_axi_rmem16_RID),
    .m00_axi_rlast(m_axi_rmem16_RLAST),
    .m00_axi_rready(m_axi_rmem16_RREADY),
    .m00_axi_rresp(m_axi_rmem16_RRESP),
    .m00_axi_rvalid(m_axi_rmem16_RVALID),
    .m00_axi_wdata(m_axi_rmem16_WDATA),
    .m00_axi_wlast(m_axi_rmem16_WLAST),
    .m00_axi_wready(m_axi_rmem16_WREADY),
    .m00_axi_wstrb(m_axi_rmem16_WSTRB),
    .m00_axi_wvalid(m_axi_rmem16_WVALID),
    .s00_axi_araddr(m_axi_rmem16___Mmap2Stream_16___mmap_ARADDR),
    .s00_axi_arburst(m_axi_rmem16___Mmap2Stream_16___mmap_ARBURST),
    .s00_axi_arcache(m_axi_rmem16___Mmap2Stream_16___mmap_ARCACHE),
    .s00_axi_arid(m_axi_rmem16___Mmap2Stream_16___mmap_ARID),
    .s00_axi_arlen(m_axi_rmem16___Mmap2Stream_16___mmap_ARLEN),
    .s00_axi_arlock(m_axi_rmem16___Mmap2Stream_16___mmap_ARLOCK),
    .s00_axi_arprot(m_axi_rmem16___Mmap2Stream_16___mmap_ARPROT),
    .s00_axi_arqos(m_axi_rmem16___Mmap2Stream_16___mmap_ARQOS),
    .s00_axi_arready(m_axi_rmem16___Mmap2Stream_16___mmap_ARREADY),
    .s00_axi_arsize(m_axi_rmem16___Mmap2Stream_16___mmap_ARSIZE),
    .s00_axi_arvalid(m_axi_rmem16___Mmap2Stream_16___mmap_ARVALID),
    .s00_axi_awaddr(m_axi_rmem16___Mmap2Stream_16___mmap_AWADDR),
    .s00_axi_awburst(m_axi_rmem16___Mmap2Stream_16___mmap_AWBURST),
    .s00_axi_awcache(m_axi_rmem16___Mmap2Stream_16___mmap_AWCACHE),
    .s00_axi_awid(m_axi_rmem16___Mmap2Stream_16___mmap_AWID),
    .s00_axi_awlen(m_axi_rmem16___Mmap2Stream_16___mmap_AWLEN),
    .s00_axi_awlock(m_axi_rmem16___Mmap2Stream_16___mmap_AWLOCK),
    .s00_axi_awprot(m_axi_rmem16___Mmap2Stream_16___mmap_AWPROT),
    .s00_axi_awqos(m_axi_rmem16___Mmap2Stream_16___mmap_AWQOS),
    .s00_axi_awready(m_axi_rmem16___Mmap2Stream_16___mmap_AWREADY),
    .s00_axi_awsize(m_axi_rmem16___Mmap2Stream_16___mmap_AWSIZE),
    .s00_axi_awvalid(m_axi_rmem16___Mmap2Stream_16___mmap_AWVALID),
    .s00_axi_bid(m_axi_rmem16___Mmap2Stream_16___mmap_BID),
    .s00_axi_bready(m_axi_rmem16___Mmap2Stream_16___mmap_BREADY),
    .s00_axi_bresp(m_axi_rmem16___Mmap2Stream_16___mmap_BRESP),
    .s00_axi_bvalid(m_axi_rmem16___Mmap2Stream_16___mmap_BVALID),
    .s00_axi_rdata(m_axi_rmem16___Mmap2Stream_16___mmap_RDATA),
    .s00_axi_rid(m_axi_rmem16___Mmap2Stream_16___mmap_RID),
    .s00_axi_rlast(m_axi_rmem16___Mmap2Stream_16___mmap_RLAST),
    .s00_axi_rready(m_axi_rmem16___Mmap2Stream_16___mmap_RREADY),
    .s00_axi_rresp(m_axi_rmem16___Mmap2Stream_16___mmap_RRESP),
    .s00_axi_rvalid(m_axi_rmem16___Mmap2Stream_16___mmap_RVALID),
    .s00_axi_wdata(m_axi_rmem16___Mmap2Stream_16___mmap_WDATA),
    .s00_axi_wlast(m_axi_rmem16___Mmap2Stream_16___mmap_WLAST),
    .s00_axi_wready(m_axi_rmem16___Mmap2Stream_16___mmap_WREADY),
    .s00_axi_wstrb(m_axi_rmem16___Mmap2Stream_16___mmap_WSTRB),
    .s00_axi_wvalid(m_axi_rmem16___Mmap2Stream_16___mmap_WVALID),
    .s01_axi_araddr(m_axi_rmem16___Stream2Mmap_16___mmap_ARADDR),
    .s01_axi_arburst(m_axi_rmem16___Stream2Mmap_16___mmap_ARBURST),
    .s01_axi_arcache(m_axi_rmem16___Stream2Mmap_16___mmap_ARCACHE),
    .s01_axi_arid(m_axi_rmem16___Stream2Mmap_16___mmap_ARID),
    .s01_axi_arlen(m_axi_rmem16___Stream2Mmap_16___mmap_ARLEN),
    .s01_axi_arlock(m_axi_rmem16___Stream2Mmap_16___mmap_ARLOCK),
    .s01_axi_arprot(m_axi_rmem16___Stream2Mmap_16___mmap_ARPROT),
    .s01_axi_arqos(m_axi_rmem16___Stream2Mmap_16___mmap_ARQOS),
    .s01_axi_arready(m_axi_rmem16___Stream2Mmap_16___mmap_ARREADY),
    .s01_axi_arsize(m_axi_rmem16___Stream2Mmap_16___mmap_ARSIZE),
    .s01_axi_arvalid(m_axi_rmem16___Stream2Mmap_16___mmap_ARVALID),
    .s01_axi_awaddr(m_axi_rmem16___Stream2Mmap_16___mmap_AWADDR),
    .s01_axi_awburst(m_axi_rmem16___Stream2Mmap_16___mmap_AWBURST),
    .s01_axi_awcache(m_axi_rmem16___Stream2Mmap_16___mmap_AWCACHE),
    .s01_axi_awid(m_axi_rmem16___Stream2Mmap_16___mmap_AWID),
    .s01_axi_awlen(m_axi_rmem16___Stream2Mmap_16___mmap_AWLEN),
    .s01_axi_awlock(m_axi_rmem16___Stream2Mmap_16___mmap_AWLOCK),
    .s01_axi_awprot(m_axi_rmem16___Stream2Mmap_16___mmap_AWPROT),
    .s01_axi_awqos(m_axi_rmem16___Stream2Mmap_16___mmap_AWQOS),
    .s01_axi_awready(m_axi_rmem16___Stream2Mmap_16___mmap_AWREADY),
    .s01_axi_awsize(m_axi_rmem16___Stream2Mmap_16___mmap_AWSIZE),
    .s01_axi_awvalid(m_axi_rmem16___Stream2Mmap_16___mmap_AWVALID),
    .s01_axi_bid(m_axi_rmem16___Stream2Mmap_16___mmap_BID),
    .s01_axi_bready(m_axi_rmem16___Stream2Mmap_16___mmap_BREADY),
    .s01_axi_bresp(m_axi_rmem16___Stream2Mmap_16___mmap_BRESP),
    .s01_axi_bvalid(m_axi_rmem16___Stream2Mmap_16___mmap_BVALID),
    .s01_axi_rdata(m_axi_rmem16___Stream2Mmap_16___mmap_RDATA),
    .s01_axi_rid(m_axi_rmem16___Stream2Mmap_16___mmap_RID),
    .s01_axi_rlast(m_axi_rmem16___Stream2Mmap_16___mmap_RLAST),
    .s01_axi_rready(m_axi_rmem16___Stream2Mmap_16___mmap_RREADY),
    .s01_axi_rresp(m_axi_rmem16___Stream2Mmap_16___mmap_RRESP),
    .s01_axi_rvalid(m_axi_rmem16___Stream2Mmap_16___mmap_RVALID),
    .s01_axi_wdata(m_axi_rmem16___Stream2Mmap_16___mmap_WDATA),
    .s01_axi_wlast(m_axi_rmem16___Stream2Mmap_16___mmap_WLAST),
    .s01_axi_wready(m_axi_rmem16___Stream2Mmap_16___mmap_WREADY),
    .s01_axi_wstrb(m_axi_rmem16___Stream2Mmap_16___mmap_WSTRB),
    .s01_axi_wvalid(m_axi_rmem16___Stream2Mmap_16___mmap_WVALID)
  );


  (* keep_hierarchy = "yes" *) axi_crossbar_2x1
  #(
    .DATA_WIDTH(512),
    .ADDR_WIDTH(64),
    .S_ID_WIDTH(1),
    .M_ID_WIDTH(2),
    .M00_ADDR_WIDTH(64),
    .M00_ISSUE(16),
    .S00_THREADS(1),
    .S01_THREADS(1)
  )
  axi_crossbar_2x1__rmem17
  (
    .clk(ap_clk),
    .rst(ap_rst_n_inv),
    .m00_axi_araddr(m_axi_rmem17_ARADDR),
    .m00_axi_arburst(m_axi_rmem17_ARBURST),
    .m00_axi_arcache(m_axi_rmem17_ARCACHE),
    .m00_axi_arid(m_axi_rmem17_ARID),
    .m00_axi_arlen(m_axi_rmem17_ARLEN),
    .m00_axi_arlock(m_axi_rmem17_ARLOCK),
    .m00_axi_arprot(m_axi_rmem17_ARPROT),
    .m00_axi_arqos(m_axi_rmem17_ARQOS),
    .m00_axi_arready(m_axi_rmem17_ARREADY),
    .m00_axi_arsize(m_axi_rmem17_ARSIZE),
    .m00_axi_arvalid(m_axi_rmem17_ARVALID),
    .m00_axi_awaddr(m_axi_rmem17_AWADDR),
    .m00_axi_awburst(m_axi_rmem17_AWBURST),
    .m00_axi_awcache(m_axi_rmem17_AWCACHE),
    .m00_axi_awid(m_axi_rmem17_AWID),
    .m00_axi_awlen(m_axi_rmem17_AWLEN),
    .m00_axi_awlock(m_axi_rmem17_AWLOCK),
    .m00_axi_awprot(m_axi_rmem17_AWPROT),
    .m00_axi_awqos(m_axi_rmem17_AWQOS),
    .m00_axi_awready(m_axi_rmem17_AWREADY),
    .m00_axi_awsize(m_axi_rmem17_AWSIZE),
    .m00_axi_awvalid(m_axi_rmem17_AWVALID),
    .m00_axi_bid(m_axi_rmem17_BID),
    .m00_axi_bready(m_axi_rmem17_BREADY),
    .m00_axi_bresp(m_axi_rmem17_BRESP),
    .m00_axi_bvalid(m_axi_rmem17_BVALID),
    .m00_axi_rdata(m_axi_rmem17_RDATA),
    .m00_axi_rid(m_axi_rmem17_RID),
    .m00_axi_rlast(m_axi_rmem17_RLAST),
    .m00_axi_rready(m_axi_rmem17_RREADY),
    .m00_axi_rresp(m_axi_rmem17_RRESP),
    .m00_axi_rvalid(m_axi_rmem17_RVALID),
    .m00_axi_wdata(m_axi_rmem17_WDATA),
    .m00_axi_wlast(m_axi_rmem17_WLAST),
    .m00_axi_wready(m_axi_rmem17_WREADY),
    .m00_axi_wstrb(m_axi_rmem17_WSTRB),
    .m00_axi_wvalid(m_axi_rmem17_WVALID),
    .s00_axi_araddr(m_axi_rmem17___Mmap2Stream_17___mmap_ARADDR),
    .s00_axi_arburst(m_axi_rmem17___Mmap2Stream_17___mmap_ARBURST),
    .s00_axi_arcache(m_axi_rmem17___Mmap2Stream_17___mmap_ARCACHE),
    .s00_axi_arid(m_axi_rmem17___Mmap2Stream_17___mmap_ARID),
    .s00_axi_arlen(m_axi_rmem17___Mmap2Stream_17___mmap_ARLEN),
    .s00_axi_arlock(m_axi_rmem17___Mmap2Stream_17___mmap_ARLOCK),
    .s00_axi_arprot(m_axi_rmem17___Mmap2Stream_17___mmap_ARPROT),
    .s00_axi_arqos(m_axi_rmem17___Mmap2Stream_17___mmap_ARQOS),
    .s00_axi_arready(m_axi_rmem17___Mmap2Stream_17___mmap_ARREADY),
    .s00_axi_arsize(m_axi_rmem17___Mmap2Stream_17___mmap_ARSIZE),
    .s00_axi_arvalid(m_axi_rmem17___Mmap2Stream_17___mmap_ARVALID),
    .s00_axi_awaddr(m_axi_rmem17___Mmap2Stream_17___mmap_AWADDR),
    .s00_axi_awburst(m_axi_rmem17___Mmap2Stream_17___mmap_AWBURST),
    .s00_axi_awcache(m_axi_rmem17___Mmap2Stream_17___mmap_AWCACHE),
    .s00_axi_awid(m_axi_rmem17___Mmap2Stream_17___mmap_AWID),
    .s00_axi_awlen(m_axi_rmem17___Mmap2Stream_17___mmap_AWLEN),
    .s00_axi_awlock(m_axi_rmem17___Mmap2Stream_17___mmap_AWLOCK),
    .s00_axi_awprot(m_axi_rmem17___Mmap2Stream_17___mmap_AWPROT),
    .s00_axi_awqos(m_axi_rmem17___Mmap2Stream_17___mmap_AWQOS),
    .s00_axi_awready(m_axi_rmem17___Mmap2Stream_17___mmap_AWREADY),
    .s00_axi_awsize(m_axi_rmem17___Mmap2Stream_17___mmap_AWSIZE),
    .s00_axi_awvalid(m_axi_rmem17___Mmap2Stream_17___mmap_AWVALID),
    .s00_axi_bid(m_axi_rmem17___Mmap2Stream_17___mmap_BID),
    .s00_axi_bready(m_axi_rmem17___Mmap2Stream_17___mmap_BREADY),
    .s00_axi_bresp(m_axi_rmem17___Mmap2Stream_17___mmap_BRESP),
    .s00_axi_bvalid(m_axi_rmem17___Mmap2Stream_17___mmap_BVALID),
    .s00_axi_rdata(m_axi_rmem17___Mmap2Stream_17___mmap_RDATA),
    .s00_axi_rid(m_axi_rmem17___Mmap2Stream_17___mmap_RID),
    .s00_axi_rlast(m_axi_rmem17___Mmap2Stream_17___mmap_RLAST),
    .s00_axi_rready(m_axi_rmem17___Mmap2Stream_17___mmap_RREADY),
    .s00_axi_rresp(m_axi_rmem17___Mmap2Stream_17___mmap_RRESP),
    .s00_axi_rvalid(m_axi_rmem17___Mmap2Stream_17___mmap_RVALID),
    .s00_axi_wdata(m_axi_rmem17___Mmap2Stream_17___mmap_WDATA),
    .s00_axi_wlast(m_axi_rmem17___Mmap2Stream_17___mmap_WLAST),
    .s00_axi_wready(m_axi_rmem17___Mmap2Stream_17___mmap_WREADY),
    .s00_axi_wstrb(m_axi_rmem17___Mmap2Stream_17___mmap_WSTRB),
    .s00_axi_wvalid(m_axi_rmem17___Mmap2Stream_17___mmap_WVALID),
    .s01_axi_araddr(m_axi_rmem17___Stream2Mmap_17___mmap_ARADDR),
    .s01_axi_arburst(m_axi_rmem17___Stream2Mmap_17___mmap_ARBURST),
    .s01_axi_arcache(m_axi_rmem17___Stream2Mmap_17___mmap_ARCACHE),
    .s01_axi_arid(m_axi_rmem17___Stream2Mmap_17___mmap_ARID),
    .s01_axi_arlen(m_axi_rmem17___Stream2Mmap_17___mmap_ARLEN),
    .s01_axi_arlock(m_axi_rmem17___Stream2Mmap_17___mmap_ARLOCK),
    .s01_axi_arprot(m_axi_rmem17___Stream2Mmap_17___mmap_ARPROT),
    .s01_axi_arqos(m_axi_rmem17___Stream2Mmap_17___mmap_ARQOS),
    .s01_axi_arready(m_axi_rmem17___Stream2Mmap_17___mmap_ARREADY),
    .s01_axi_arsize(m_axi_rmem17___Stream2Mmap_17___mmap_ARSIZE),
    .s01_axi_arvalid(m_axi_rmem17___Stream2Mmap_17___mmap_ARVALID),
    .s01_axi_awaddr(m_axi_rmem17___Stream2Mmap_17___mmap_AWADDR),
    .s01_axi_awburst(m_axi_rmem17___Stream2Mmap_17___mmap_AWBURST),
    .s01_axi_awcache(m_axi_rmem17___Stream2Mmap_17___mmap_AWCACHE),
    .s01_axi_awid(m_axi_rmem17___Stream2Mmap_17___mmap_AWID),
    .s01_axi_awlen(m_axi_rmem17___Stream2Mmap_17___mmap_AWLEN),
    .s01_axi_awlock(m_axi_rmem17___Stream2Mmap_17___mmap_AWLOCK),
    .s01_axi_awprot(m_axi_rmem17___Stream2Mmap_17___mmap_AWPROT),
    .s01_axi_awqos(m_axi_rmem17___Stream2Mmap_17___mmap_AWQOS),
    .s01_axi_awready(m_axi_rmem17___Stream2Mmap_17___mmap_AWREADY),
    .s01_axi_awsize(m_axi_rmem17___Stream2Mmap_17___mmap_AWSIZE),
    .s01_axi_awvalid(m_axi_rmem17___Stream2Mmap_17___mmap_AWVALID),
    .s01_axi_bid(m_axi_rmem17___Stream2Mmap_17___mmap_BID),
    .s01_axi_bready(m_axi_rmem17___Stream2Mmap_17___mmap_BREADY),
    .s01_axi_bresp(m_axi_rmem17___Stream2Mmap_17___mmap_BRESP),
    .s01_axi_bvalid(m_axi_rmem17___Stream2Mmap_17___mmap_BVALID),
    .s01_axi_rdata(m_axi_rmem17___Stream2Mmap_17___mmap_RDATA),
    .s01_axi_rid(m_axi_rmem17___Stream2Mmap_17___mmap_RID),
    .s01_axi_rlast(m_axi_rmem17___Stream2Mmap_17___mmap_RLAST),
    .s01_axi_rready(m_axi_rmem17___Stream2Mmap_17___mmap_RREADY),
    .s01_axi_rresp(m_axi_rmem17___Stream2Mmap_17___mmap_RRESP),
    .s01_axi_rvalid(m_axi_rmem17___Stream2Mmap_17___mmap_RVALID),
    .s01_axi_wdata(m_axi_rmem17___Stream2Mmap_17___mmap_WDATA),
    .s01_axi_wlast(m_axi_rmem17___Stream2Mmap_17___mmap_WLAST),
    .s01_axi_wready(m_axi_rmem17___Stream2Mmap_17___mmap_WREADY),
    .s01_axi_wstrb(m_axi_rmem17___Stream2Mmap_17___mmap_WSTRB),
    .s01_axi_wvalid(m_axi_rmem17___Stream2Mmap_17___mmap_WVALID)
  );


  (* keep_hierarchy = "yes" *) axi_crossbar_2x1
  #(
    .DATA_WIDTH(512),
    .ADDR_WIDTH(64),
    .S_ID_WIDTH(1),
    .M_ID_WIDTH(2),
    .M00_ADDR_WIDTH(64),
    .M00_ISSUE(16),
    .S00_THREADS(1),
    .S01_THREADS(1)
  )
  axi_crossbar_2x1__rmem18
  (
    .clk(ap_clk),
    .rst(ap_rst_n_inv),
    .m00_axi_araddr(m_axi_rmem18_ARADDR),
    .m00_axi_arburst(m_axi_rmem18_ARBURST),
    .m00_axi_arcache(m_axi_rmem18_ARCACHE),
    .m00_axi_arid(m_axi_rmem18_ARID),
    .m00_axi_arlen(m_axi_rmem18_ARLEN),
    .m00_axi_arlock(m_axi_rmem18_ARLOCK),
    .m00_axi_arprot(m_axi_rmem18_ARPROT),
    .m00_axi_arqos(m_axi_rmem18_ARQOS),
    .m00_axi_arready(m_axi_rmem18_ARREADY),
    .m00_axi_arsize(m_axi_rmem18_ARSIZE),
    .m00_axi_arvalid(m_axi_rmem18_ARVALID),
    .m00_axi_awaddr(m_axi_rmem18_AWADDR),
    .m00_axi_awburst(m_axi_rmem18_AWBURST),
    .m00_axi_awcache(m_axi_rmem18_AWCACHE),
    .m00_axi_awid(m_axi_rmem18_AWID),
    .m00_axi_awlen(m_axi_rmem18_AWLEN),
    .m00_axi_awlock(m_axi_rmem18_AWLOCK),
    .m00_axi_awprot(m_axi_rmem18_AWPROT),
    .m00_axi_awqos(m_axi_rmem18_AWQOS),
    .m00_axi_awready(m_axi_rmem18_AWREADY),
    .m00_axi_awsize(m_axi_rmem18_AWSIZE),
    .m00_axi_awvalid(m_axi_rmem18_AWVALID),
    .m00_axi_bid(m_axi_rmem18_BID),
    .m00_axi_bready(m_axi_rmem18_BREADY),
    .m00_axi_bresp(m_axi_rmem18_BRESP),
    .m00_axi_bvalid(m_axi_rmem18_BVALID),
    .m00_axi_rdata(m_axi_rmem18_RDATA),
    .m00_axi_rid(m_axi_rmem18_RID),
    .m00_axi_rlast(m_axi_rmem18_RLAST),
    .m00_axi_rready(m_axi_rmem18_RREADY),
    .m00_axi_rresp(m_axi_rmem18_RRESP),
    .m00_axi_rvalid(m_axi_rmem18_RVALID),
    .m00_axi_wdata(m_axi_rmem18_WDATA),
    .m00_axi_wlast(m_axi_rmem18_WLAST),
    .m00_axi_wready(m_axi_rmem18_WREADY),
    .m00_axi_wstrb(m_axi_rmem18_WSTRB),
    .m00_axi_wvalid(m_axi_rmem18_WVALID),
    .s00_axi_araddr(m_axi_rmem18___Mmap2Stream_18___mmap_ARADDR),
    .s00_axi_arburst(m_axi_rmem18___Mmap2Stream_18___mmap_ARBURST),
    .s00_axi_arcache(m_axi_rmem18___Mmap2Stream_18___mmap_ARCACHE),
    .s00_axi_arid(m_axi_rmem18___Mmap2Stream_18___mmap_ARID),
    .s00_axi_arlen(m_axi_rmem18___Mmap2Stream_18___mmap_ARLEN),
    .s00_axi_arlock(m_axi_rmem18___Mmap2Stream_18___mmap_ARLOCK),
    .s00_axi_arprot(m_axi_rmem18___Mmap2Stream_18___mmap_ARPROT),
    .s00_axi_arqos(m_axi_rmem18___Mmap2Stream_18___mmap_ARQOS),
    .s00_axi_arready(m_axi_rmem18___Mmap2Stream_18___mmap_ARREADY),
    .s00_axi_arsize(m_axi_rmem18___Mmap2Stream_18___mmap_ARSIZE),
    .s00_axi_arvalid(m_axi_rmem18___Mmap2Stream_18___mmap_ARVALID),
    .s00_axi_awaddr(m_axi_rmem18___Mmap2Stream_18___mmap_AWADDR),
    .s00_axi_awburst(m_axi_rmem18___Mmap2Stream_18___mmap_AWBURST),
    .s00_axi_awcache(m_axi_rmem18___Mmap2Stream_18___mmap_AWCACHE),
    .s00_axi_awid(m_axi_rmem18___Mmap2Stream_18___mmap_AWID),
    .s00_axi_awlen(m_axi_rmem18___Mmap2Stream_18___mmap_AWLEN),
    .s00_axi_awlock(m_axi_rmem18___Mmap2Stream_18___mmap_AWLOCK),
    .s00_axi_awprot(m_axi_rmem18___Mmap2Stream_18___mmap_AWPROT),
    .s00_axi_awqos(m_axi_rmem18___Mmap2Stream_18___mmap_AWQOS),
    .s00_axi_awready(m_axi_rmem18___Mmap2Stream_18___mmap_AWREADY),
    .s00_axi_awsize(m_axi_rmem18___Mmap2Stream_18___mmap_AWSIZE),
    .s00_axi_awvalid(m_axi_rmem18___Mmap2Stream_18___mmap_AWVALID),
    .s00_axi_bid(m_axi_rmem18___Mmap2Stream_18___mmap_BID),
    .s00_axi_bready(m_axi_rmem18___Mmap2Stream_18___mmap_BREADY),
    .s00_axi_bresp(m_axi_rmem18___Mmap2Stream_18___mmap_BRESP),
    .s00_axi_bvalid(m_axi_rmem18___Mmap2Stream_18___mmap_BVALID),
    .s00_axi_rdata(m_axi_rmem18___Mmap2Stream_18___mmap_RDATA),
    .s00_axi_rid(m_axi_rmem18___Mmap2Stream_18___mmap_RID),
    .s00_axi_rlast(m_axi_rmem18___Mmap2Stream_18___mmap_RLAST),
    .s00_axi_rready(m_axi_rmem18___Mmap2Stream_18___mmap_RREADY),
    .s00_axi_rresp(m_axi_rmem18___Mmap2Stream_18___mmap_RRESP),
    .s00_axi_rvalid(m_axi_rmem18___Mmap2Stream_18___mmap_RVALID),
    .s00_axi_wdata(m_axi_rmem18___Mmap2Stream_18___mmap_WDATA),
    .s00_axi_wlast(m_axi_rmem18___Mmap2Stream_18___mmap_WLAST),
    .s00_axi_wready(m_axi_rmem18___Mmap2Stream_18___mmap_WREADY),
    .s00_axi_wstrb(m_axi_rmem18___Mmap2Stream_18___mmap_WSTRB),
    .s00_axi_wvalid(m_axi_rmem18___Mmap2Stream_18___mmap_WVALID),
    .s01_axi_araddr(m_axi_rmem18___Stream2Mmap_18___mmap_ARADDR),
    .s01_axi_arburst(m_axi_rmem18___Stream2Mmap_18___mmap_ARBURST),
    .s01_axi_arcache(m_axi_rmem18___Stream2Mmap_18___mmap_ARCACHE),
    .s01_axi_arid(m_axi_rmem18___Stream2Mmap_18___mmap_ARID),
    .s01_axi_arlen(m_axi_rmem18___Stream2Mmap_18___mmap_ARLEN),
    .s01_axi_arlock(m_axi_rmem18___Stream2Mmap_18___mmap_ARLOCK),
    .s01_axi_arprot(m_axi_rmem18___Stream2Mmap_18___mmap_ARPROT),
    .s01_axi_arqos(m_axi_rmem18___Stream2Mmap_18___mmap_ARQOS),
    .s01_axi_arready(m_axi_rmem18___Stream2Mmap_18___mmap_ARREADY),
    .s01_axi_arsize(m_axi_rmem18___Stream2Mmap_18___mmap_ARSIZE),
    .s01_axi_arvalid(m_axi_rmem18___Stream2Mmap_18___mmap_ARVALID),
    .s01_axi_awaddr(m_axi_rmem18___Stream2Mmap_18___mmap_AWADDR),
    .s01_axi_awburst(m_axi_rmem18___Stream2Mmap_18___mmap_AWBURST),
    .s01_axi_awcache(m_axi_rmem18___Stream2Mmap_18___mmap_AWCACHE),
    .s01_axi_awid(m_axi_rmem18___Stream2Mmap_18___mmap_AWID),
    .s01_axi_awlen(m_axi_rmem18___Stream2Mmap_18___mmap_AWLEN),
    .s01_axi_awlock(m_axi_rmem18___Stream2Mmap_18___mmap_AWLOCK),
    .s01_axi_awprot(m_axi_rmem18___Stream2Mmap_18___mmap_AWPROT),
    .s01_axi_awqos(m_axi_rmem18___Stream2Mmap_18___mmap_AWQOS),
    .s01_axi_awready(m_axi_rmem18___Stream2Mmap_18___mmap_AWREADY),
    .s01_axi_awsize(m_axi_rmem18___Stream2Mmap_18___mmap_AWSIZE),
    .s01_axi_awvalid(m_axi_rmem18___Stream2Mmap_18___mmap_AWVALID),
    .s01_axi_bid(m_axi_rmem18___Stream2Mmap_18___mmap_BID),
    .s01_axi_bready(m_axi_rmem18___Stream2Mmap_18___mmap_BREADY),
    .s01_axi_bresp(m_axi_rmem18___Stream2Mmap_18___mmap_BRESP),
    .s01_axi_bvalid(m_axi_rmem18___Stream2Mmap_18___mmap_BVALID),
    .s01_axi_rdata(m_axi_rmem18___Stream2Mmap_18___mmap_RDATA),
    .s01_axi_rid(m_axi_rmem18___Stream2Mmap_18___mmap_RID),
    .s01_axi_rlast(m_axi_rmem18___Stream2Mmap_18___mmap_RLAST),
    .s01_axi_rready(m_axi_rmem18___Stream2Mmap_18___mmap_RREADY),
    .s01_axi_rresp(m_axi_rmem18___Stream2Mmap_18___mmap_RRESP),
    .s01_axi_rvalid(m_axi_rmem18___Stream2Mmap_18___mmap_RVALID),
    .s01_axi_wdata(m_axi_rmem18___Stream2Mmap_18___mmap_WDATA),
    .s01_axi_wlast(m_axi_rmem18___Stream2Mmap_18___mmap_WLAST),
    .s01_axi_wready(m_axi_rmem18___Stream2Mmap_18___mmap_WREADY),
    .s01_axi_wstrb(m_axi_rmem18___Stream2Mmap_18___mmap_WSTRB),
    .s01_axi_wvalid(m_axi_rmem18___Stream2Mmap_18___mmap_WVALID)
  );


  (* keep_hierarchy = "yes" *) axi_crossbar_2x1
  #(
    .DATA_WIDTH(512),
    .ADDR_WIDTH(64),
    .S_ID_WIDTH(1),
    .M_ID_WIDTH(2),
    .M00_ADDR_WIDTH(64),
    .M00_ISSUE(16),
    .S00_THREADS(1),
    .S01_THREADS(1)
  )
  axi_crossbar_2x1__rmem19
  (
    .clk(ap_clk),
    .rst(ap_rst_n_inv),
    .m00_axi_araddr(m_axi_rmem19_ARADDR),
    .m00_axi_arburst(m_axi_rmem19_ARBURST),
    .m00_axi_arcache(m_axi_rmem19_ARCACHE),
    .m00_axi_arid(m_axi_rmem19_ARID),
    .m00_axi_arlen(m_axi_rmem19_ARLEN),
    .m00_axi_arlock(m_axi_rmem19_ARLOCK),
    .m00_axi_arprot(m_axi_rmem19_ARPROT),
    .m00_axi_arqos(m_axi_rmem19_ARQOS),
    .m00_axi_arready(m_axi_rmem19_ARREADY),
    .m00_axi_arsize(m_axi_rmem19_ARSIZE),
    .m00_axi_arvalid(m_axi_rmem19_ARVALID),
    .m00_axi_awaddr(m_axi_rmem19_AWADDR),
    .m00_axi_awburst(m_axi_rmem19_AWBURST),
    .m00_axi_awcache(m_axi_rmem19_AWCACHE),
    .m00_axi_awid(m_axi_rmem19_AWID),
    .m00_axi_awlen(m_axi_rmem19_AWLEN),
    .m00_axi_awlock(m_axi_rmem19_AWLOCK),
    .m00_axi_awprot(m_axi_rmem19_AWPROT),
    .m00_axi_awqos(m_axi_rmem19_AWQOS),
    .m00_axi_awready(m_axi_rmem19_AWREADY),
    .m00_axi_awsize(m_axi_rmem19_AWSIZE),
    .m00_axi_awvalid(m_axi_rmem19_AWVALID),
    .m00_axi_bid(m_axi_rmem19_BID),
    .m00_axi_bready(m_axi_rmem19_BREADY),
    .m00_axi_bresp(m_axi_rmem19_BRESP),
    .m00_axi_bvalid(m_axi_rmem19_BVALID),
    .m00_axi_rdata(m_axi_rmem19_RDATA),
    .m00_axi_rid(m_axi_rmem19_RID),
    .m00_axi_rlast(m_axi_rmem19_RLAST),
    .m00_axi_rready(m_axi_rmem19_RREADY),
    .m00_axi_rresp(m_axi_rmem19_RRESP),
    .m00_axi_rvalid(m_axi_rmem19_RVALID),
    .m00_axi_wdata(m_axi_rmem19_WDATA),
    .m00_axi_wlast(m_axi_rmem19_WLAST),
    .m00_axi_wready(m_axi_rmem19_WREADY),
    .m00_axi_wstrb(m_axi_rmem19_WSTRB),
    .m00_axi_wvalid(m_axi_rmem19_WVALID),
    .s00_axi_araddr(m_axi_rmem19___Mmap2Stream_19___mmap_ARADDR),
    .s00_axi_arburst(m_axi_rmem19___Mmap2Stream_19___mmap_ARBURST),
    .s00_axi_arcache(m_axi_rmem19___Mmap2Stream_19___mmap_ARCACHE),
    .s00_axi_arid(m_axi_rmem19___Mmap2Stream_19___mmap_ARID),
    .s00_axi_arlen(m_axi_rmem19___Mmap2Stream_19___mmap_ARLEN),
    .s00_axi_arlock(m_axi_rmem19___Mmap2Stream_19___mmap_ARLOCK),
    .s00_axi_arprot(m_axi_rmem19___Mmap2Stream_19___mmap_ARPROT),
    .s00_axi_arqos(m_axi_rmem19___Mmap2Stream_19___mmap_ARQOS),
    .s00_axi_arready(m_axi_rmem19___Mmap2Stream_19___mmap_ARREADY),
    .s00_axi_arsize(m_axi_rmem19___Mmap2Stream_19___mmap_ARSIZE),
    .s00_axi_arvalid(m_axi_rmem19___Mmap2Stream_19___mmap_ARVALID),
    .s00_axi_awaddr(m_axi_rmem19___Mmap2Stream_19___mmap_AWADDR),
    .s00_axi_awburst(m_axi_rmem19___Mmap2Stream_19___mmap_AWBURST),
    .s00_axi_awcache(m_axi_rmem19___Mmap2Stream_19___mmap_AWCACHE),
    .s00_axi_awid(m_axi_rmem19___Mmap2Stream_19___mmap_AWID),
    .s00_axi_awlen(m_axi_rmem19___Mmap2Stream_19___mmap_AWLEN),
    .s00_axi_awlock(m_axi_rmem19___Mmap2Stream_19___mmap_AWLOCK),
    .s00_axi_awprot(m_axi_rmem19___Mmap2Stream_19___mmap_AWPROT),
    .s00_axi_awqos(m_axi_rmem19___Mmap2Stream_19___mmap_AWQOS),
    .s00_axi_awready(m_axi_rmem19___Mmap2Stream_19___mmap_AWREADY),
    .s00_axi_awsize(m_axi_rmem19___Mmap2Stream_19___mmap_AWSIZE),
    .s00_axi_awvalid(m_axi_rmem19___Mmap2Stream_19___mmap_AWVALID),
    .s00_axi_bid(m_axi_rmem19___Mmap2Stream_19___mmap_BID),
    .s00_axi_bready(m_axi_rmem19___Mmap2Stream_19___mmap_BREADY),
    .s00_axi_bresp(m_axi_rmem19___Mmap2Stream_19___mmap_BRESP),
    .s00_axi_bvalid(m_axi_rmem19___Mmap2Stream_19___mmap_BVALID),
    .s00_axi_rdata(m_axi_rmem19___Mmap2Stream_19___mmap_RDATA),
    .s00_axi_rid(m_axi_rmem19___Mmap2Stream_19___mmap_RID),
    .s00_axi_rlast(m_axi_rmem19___Mmap2Stream_19___mmap_RLAST),
    .s00_axi_rready(m_axi_rmem19___Mmap2Stream_19___mmap_RREADY),
    .s00_axi_rresp(m_axi_rmem19___Mmap2Stream_19___mmap_RRESP),
    .s00_axi_rvalid(m_axi_rmem19___Mmap2Stream_19___mmap_RVALID),
    .s00_axi_wdata(m_axi_rmem19___Mmap2Stream_19___mmap_WDATA),
    .s00_axi_wlast(m_axi_rmem19___Mmap2Stream_19___mmap_WLAST),
    .s00_axi_wready(m_axi_rmem19___Mmap2Stream_19___mmap_WREADY),
    .s00_axi_wstrb(m_axi_rmem19___Mmap2Stream_19___mmap_WSTRB),
    .s00_axi_wvalid(m_axi_rmem19___Mmap2Stream_19___mmap_WVALID),
    .s01_axi_araddr(m_axi_rmem19___Stream2Mmap_19___mmap_ARADDR),
    .s01_axi_arburst(m_axi_rmem19___Stream2Mmap_19___mmap_ARBURST),
    .s01_axi_arcache(m_axi_rmem19___Stream2Mmap_19___mmap_ARCACHE),
    .s01_axi_arid(m_axi_rmem19___Stream2Mmap_19___mmap_ARID),
    .s01_axi_arlen(m_axi_rmem19___Stream2Mmap_19___mmap_ARLEN),
    .s01_axi_arlock(m_axi_rmem19___Stream2Mmap_19___mmap_ARLOCK),
    .s01_axi_arprot(m_axi_rmem19___Stream2Mmap_19___mmap_ARPROT),
    .s01_axi_arqos(m_axi_rmem19___Stream2Mmap_19___mmap_ARQOS),
    .s01_axi_arready(m_axi_rmem19___Stream2Mmap_19___mmap_ARREADY),
    .s01_axi_arsize(m_axi_rmem19___Stream2Mmap_19___mmap_ARSIZE),
    .s01_axi_arvalid(m_axi_rmem19___Stream2Mmap_19___mmap_ARVALID),
    .s01_axi_awaddr(m_axi_rmem19___Stream2Mmap_19___mmap_AWADDR),
    .s01_axi_awburst(m_axi_rmem19___Stream2Mmap_19___mmap_AWBURST),
    .s01_axi_awcache(m_axi_rmem19___Stream2Mmap_19___mmap_AWCACHE),
    .s01_axi_awid(m_axi_rmem19___Stream2Mmap_19___mmap_AWID),
    .s01_axi_awlen(m_axi_rmem19___Stream2Mmap_19___mmap_AWLEN),
    .s01_axi_awlock(m_axi_rmem19___Stream2Mmap_19___mmap_AWLOCK),
    .s01_axi_awprot(m_axi_rmem19___Stream2Mmap_19___mmap_AWPROT),
    .s01_axi_awqos(m_axi_rmem19___Stream2Mmap_19___mmap_AWQOS),
    .s01_axi_awready(m_axi_rmem19___Stream2Mmap_19___mmap_AWREADY),
    .s01_axi_awsize(m_axi_rmem19___Stream2Mmap_19___mmap_AWSIZE),
    .s01_axi_awvalid(m_axi_rmem19___Stream2Mmap_19___mmap_AWVALID),
    .s01_axi_bid(m_axi_rmem19___Stream2Mmap_19___mmap_BID),
    .s01_axi_bready(m_axi_rmem19___Stream2Mmap_19___mmap_BREADY),
    .s01_axi_bresp(m_axi_rmem19___Stream2Mmap_19___mmap_BRESP),
    .s01_axi_bvalid(m_axi_rmem19___Stream2Mmap_19___mmap_BVALID),
    .s01_axi_rdata(m_axi_rmem19___Stream2Mmap_19___mmap_RDATA),
    .s01_axi_rid(m_axi_rmem19___Stream2Mmap_19___mmap_RID),
    .s01_axi_rlast(m_axi_rmem19___Stream2Mmap_19___mmap_RLAST),
    .s01_axi_rready(m_axi_rmem19___Stream2Mmap_19___mmap_RREADY),
    .s01_axi_rresp(m_axi_rmem19___Stream2Mmap_19___mmap_RRESP),
    .s01_axi_rvalid(m_axi_rmem19___Stream2Mmap_19___mmap_RVALID),
    .s01_axi_wdata(m_axi_rmem19___Stream2Mmap_19___mmap_WDATA),
    .s01_axi_wlast(m_axi_rmem19___Stream2Mmap_19___mmap_WLAST),
    .s01_axi_wready(m_axi_rmem19___Stream2Mmap_19___mmap_WREADY),
    .s01_axi_wstrb(m_axi_rmem19___Stream2Mmap_19___mmap_WSTRB),
    .s01_axi_wvalid(m_axi_rmem19___Stream2Mmap_19___mmap_WVALID)
  );


  (* keep_hierarchy = "yes" *) axi_crossbar_2x1
  #(
    .DATA_WIDTH(512),
    .ADDR_WIDTH(64),
    .S_ID_WIDTH(1),
    .M_ID_WIDTH(2),
    .M00_ADDR_WIDTH(64),
    .M00_ISSUE(16),
    .S00_THREADS(1),
    .S01_THREADS(1)
  )
  axi_crossbar_2x1__rmem20
  (
    .clk(ap_clk),
    .rst(ap_rst_n_inv),
    .m00_axi_araddr(m_axi_rmem20_ARADDR),
    .m00_axi_arburst(m_axi_rmem20_ARBURST),
    .m00_axi_arcache(m_axi_rmem20_ARCACHE),
    .m00_axi_arid(m_axi_rmem20_ARID),
    .m00_axi_arlen(m_axi_rmem20_ARLEN),
    .m00_axi_arlock(m_axi_rmem20_ARLOCK),
    .m00_axi_arprot(m_axi_rmem20_ARPROT),
    .m00_axi_arqos(m_axi_rmem20_ARQOS),
    .m00_axi_arready(m_axi_rmem20_ARREADY),
    .m00_axi_arsize(m_axi_rmem20_ARSIZE),
    .m00_axi_arvalid(m_axi_rmem20_ARVALID),
    .m00_axi_awaddr(m_axi_rmem20_AWADDR),
    .m00_axi_awburst(m_axi_rmem20_AWBURST),
    .m00_axi_awcache(m_axi_rmem20_AWCACHE),
    .m00_axi_awid(m_axi_rmem20_AWID),
    .m00_axi_awlen(m_axi_rmem20_AWLEN),
    .m00_axi_awlock(m_axi_rmem20_AWLOCK),
    .m00_axi_awprot(m_axi_rmem20_AWPROT),
    .m00_axi_awqos(m_axi_rmem20_AWQOS),
    .m00_axi_awready(m_axi_rmem20_AWREADY),
    .m00_axi_awsize(m_axi_rmem20_AWSIZE),
    .m00_axi_awvalid(m_axi_rmem20_AWVALID),
    .m00_axi_bid(m_axi_rmem20_BID),
    .m00_axi_bready(m_axi_rmem20_BREADY),
    .m00_axi_bresp(m_axi_rmem20_BRESP),
    .m00_axi_bvalid(m_axi_rmem20_BVALID),
    .m00_axi_rdata(m_axi_rmem20_RDATA),
    .m00_axi_rid(m_axi_rmem20_RID),
    .m00_axi_rlast(m_axi_rmem20_RLAST),
    .m00_axi_rready(m_axi_rmem20_RREADY),
    .m00_axi_rresp(m_axi_rmem20_RRESP),
    .m00_axi_rvalid(m_axi_rmem20_RVALID),
    .m00_axi_wdata(m_axi_rmem20_WDATA),
    .m00_axi_wlast(m_axi_rmem20_WLAST),
    .m00_axi_wready(m_axi_rmem20_WREADY),
    .m00_axi_wstrb(m_axi_rmem20_WSTRB),
    .m00_axi_wvalid(m_axi_rmem20_WVALID),
    .s00_axi_araddr(m_axi_rmem20___Mmap2Stream_20___mmap_ARADDR),
    .s00_axi_arburst(m_axi_rmem20___Mmap2Stream_20___mmap_ARBURST),
    .s00_axi_arcache(m_axi_rmem20___Mmap2Stream_20___mmap_ARCACHE),
    .s00_axi_arid(m_axi_rmem20___Mmap2Stream_20___mmap_ARID),
    .s00_axi_arlen(m_axi_rmem20___Mmap2Stream_20___mmap_ARLEN),
    .s00_axi_arlock(m_axi_rmem20___Mmap2Stream_20___mmap_ARLOCK),
    .s00_axi_arprot(m_axi_rmem20___Mmap2Stream_20___mmap_ARPROT),
    .s00_axi_arqos(m_axi_rmem20___Mmap2Stream_20___mmap_ARQOS),
    .s00_axi_arready(m_axi_rmem20___Mmap2Stream_20___mmap_ARREADY),
    .s00_axi_arsize(m_axi_rmem20___Mmap2Stream_20___mmap_ARSIZE),
    .s00_axi_arvalid(m_axi_rmem20___Mmap2Stream_20___mmap_ARVALID),
    .s00_axi_awaddr(m_axi_rmem20___Mmap2Stream_20___mmap_AWADDR),
    .s00_axi_awburst(m_axi_rmem20___Mmap2Stream_20___mmap_AWBURST),
    .s00_axi_awcache(m_axi_rmem20___Mmap2Stream_20___mmap_AWCACHE),
    .s00_axi_awid(m_axi_rmem20___Mmap2Stream_20___mmap_AWID),
    .s00_axi_awlen(m_axi_rmem20___Mmap2Stream_20___mmap_AWLEN),
    .s00_axi_awlock(m_axi_rmem20___Mmap2Stream_20___mmap_AWLOCK),
    .s00_axi_awprot(m_axi_rmem20___Mmap2Stream_20___mmap_AWPROT),
    .s00_axi_awqos(m_axi_rmem20___Mmap2Stream_20___mmap_AWQOS),
    .s00_axi_awready(m_axi_rmem20___Mmap2Stream_20___mmap_AWREADY),
    .s00_axi_awsize(m_axi_rmem20___Mmap2Stream_20___mmap_AWSIZE),
    .s00_axi_awvalid(m_axi_rmem20___Mmap2Stream_20___mmap_AWVALID),
    .s00_axi_bid(m_axi_rmem20___Mmap2Stream_20___mmap_BID),
    .s00_axi_bready(m_axi_rmem20___Mmap2Stream_20___mmap_BREADY),
    .s00_axi_bresp(m_axi_rmem20___Mmap2Stream_20___mmap_BRESP),
    .s00_axi_bvalid(m_axi_rmem20___Mmap2Stream_20___mmap_BVALID),
    .s00_axi_rdata(m_axi_rmem20___Mmap2Stream_20___mmap_RDATA),
    .s00_axi_rid(m_axi_rmem20___Mmap2Stream_20___mmap_RID),
    .s00_axi_rlast(m_axi_rmem20___Mmap2Stream_20___mmap_RLAST),
    .s00_axi_rready(m_axi_rmem20___Mmap2Stream_20___mmap_RREADY),
    .s00_axi_rresp(m_axi_rmem20___Mmap2Stream_20___mmap_RRESP),
    .s00_axi_rvalid(m_axi_rmem20___Mmap2Stream_20___mmap_RVALID),
    .s00_axi_wdata(m_axi_rmem20___Mmap2Stream_20___mmap_WDATA),
    .s00_axi_wlast(m_axi_rmem20___Mmap2Stream_20___mmap_WLAST),
    .s00_axi_wready(m_axi_rmem20___Mmap2Stream_20___mmap_WREADY),
    .s00_axi_wstrb(m_axi_rmem20___Mmap2Stream_20___mmap_WSTRB),
    .s00_axi_wvalid(m_axi_rmem20___Mmap2Stream_20___mmap_WVALID),
    .s01_axi_araddr(m_axi_rmem20___Stream2Mmap_20___mmap_ARADDR),
    .s01_axi_arburst(m_axi_rmem20___Stream2Mmap_20___mmap_ARBURST),
    .s01_axi_arcache(m_axi_rmem20___Stream2Mmap_20___mmap_ARCACHE),
    .s01_axi_arid(m_axi_rmem20___Stream2Mmap_20___mmap_ARID),
    .s01_axi_arlen(m_axi_rmem20___Stream2Mmap_20___mmap_ARLEN),
    .s01_axi_arlock(m_axi_rmem20___Stream2Mmap_20___mmap_ARLOCK),
    .s01_axi_arprot(m_axi_rmem20___Stream2Mmap_20___mmap_ARPROT),
    .s01_axi_arqos(m_axi_rmem20___Stream2Mmap_20___mmap_ARQOS),
    .s01_axi_arready(m_axi_rmem20___Stream2Mmap_20___mmap_ARREADY),
    .s01_axi_arsize(m_axi_rmem20___Stream2Mmap_20___mmap_ARSIZE),
    .s01_axi_arvalid(m_axi_rmem20___Stream2Mmap_20___mmap_ARVALID),
    .s01_axi_awaddr(m_axi_rmem20___Stream2Mmap_20___mmap_AWADDR),
    .s01_axi_awburst(m_axi_rmem20___Stream2Mmap_20___mmap_AWBURST),
    .s01_axi_awcache(m_axi_rmem20___Stream2Mmap_20___mmap_AWCACHE),
    .s01_axi_awid(m_axi_rmem20___Stream2Mmap_20___mmap_AWID),
    .s01_axi_awlen(m_axi_rmem20___Stream2Mmap_20___mmap_AWLEN),
    .s01_axi_awlock(m_axi_rmem20___Stream2Mmap_20___mmap_AWLOCK),
    .s01_axi_awprot(m_axi_rmem20___Stream2Mmap_20___mmap_AWPROT),
    .s01_axi_awqos(m_axi_rmem20___Stream2Mmap_20___mmap_AWQOS),
    .s01_axi_awready(m_axi_rmem20___Stream2Mmap_20___mmap_AWREADY),
    .s01_axi_awsize(m_axi_rmem20___Stream2Mmap_20___mmap_AWSIZE),
    .s01_axi_awvalid(m_axi_rmem20___Stream2Mmap_20___mmap_AWVALID),
    .s01_axi_bid(m_axi_rmem20___Stream2Mmap_20___mmap_BID),
    .s01_axi_bready(m_axi_rmem20___Stream2Mmap_20___mmap_BREADY),
    .s01_axi_bresp(m_axi_rmem20___Stream2Mmap_20___mmap_BRESP),
    .s01_axi_bvalid(m_axi_rmem20___Stream2Mmap_20___mmap_BVALID),
    .s01_axi_rdata(m_axi_rmem20___Stream2Mmap_20___mmap_RDATA),
    .s01_axi_rid(m_axi_rmem20___Stream2Mmap_20___mmap_RID),
    .s01_axi_rlast(m_axi_rmem20___Stream2Mmap_20___mmap_RLAST),
    .s01_axi_rready(m_axi_rmem20___Stream2Mmap_20___mmap_RREADY),
    .s01_axi_rresp(m_axi_rmem20___Stream2Mmap_20___mmap_RRESP),
    .s01_axi_rvalid(m_axi_rmem20___Stream2Mmap_20___mmap_RVALID),
    .s01_axi_wdata(m_axi_rmem20___Stream2Mmap_20___mmap_WDATA),
    .s01_axi_wlast(m_axi_rmem20___Stream2Mmap_20___mmap_WLAST),
    .s01_axi_wready(m_axi_rmem20___Stream2Mmap_20___mmap_WREADY),
    .s01_axi_wstrb(m_axi_rmem20___Stream2Mmap_20___mmap_WSTRB),
    .s01_axi_wvalid(m_axi_rmem20___Stream2Mmap_20___mmap_WVALID)
  );


  (* keep_hierarchy = "yes" *) axi_crossbar_2x1
  #(
    .DATA_WIDTH(512),
    .ADDR_WIDTH(64),
    .S_ID_WIDTH(1),
    .M_ID_WIDTH(2),
    .M00_ADDR_WIDTH(64),
    .M00_ISSUE(16),
    .S00_THREADS(1),
    .S01_THREADS(1)
  )
  axi_crossbar_2x1__rmem21
  (
    .clk(ap_clk),
    .rst(ap_rst_n_inv),
    .m00_axi_araddr(m_axi_rmem21_ARADDR),
    .m00_axi_arburst(m_axi_rmem21_ARBURST),
    .m00_axi_arcache(m_axi_rmem21_ARCACHE),
    .m00_axi_arid(m_axi_rmem21_ARID),
    .m00_axi_arlen(m_axi_rmem21_ARLEN),
    .m00_axi_arlock(m_axi_rmem21_ARLOCK),
    .m00_axi_arprot(m_axi_rmem21_ARPROT),
    .m00_axi_arqos(m_axi_rmem21_ARQOS),
    .m00_axi_arready(m_axi_rmem21_ARREADY),
    .m00_axi_arsize(m_axi_rmem21_ARSIZE),
    .m00_axi_arvalid(m_axi_rmem21_ARVALID),
    .m00_axi_awaddr(m_axi_rmem21_AWADDR),
    .m00_axi_awburst(m_axi_rmem21_AWBURST),
    .m00_axi_awcache(m_axi_rmem21_AWCACHE),
    .m00_axi_awid(m_axi_rmem21_AWID),
    .m00_axi_awlen(m_axi_rmem21_AWLEN),
    .m00_axi_awlock(m_axi_rmem21_AWLOCK),
    .m00_axi_awprot(m_axi_rmem21_AWPROT),
    .m00_axi_awqos(m_axi_rmem21_AWQOS),
    .m00_axi_awready(m_axi_rmem21_AWREADY),
    .m00_axi_awsize(m_axi_rmem21_AWSIZE),
    .m00_axi_awvalid(m_axi_rmem21_AWVALID),
    .m00_axi_bid(m_axi_rmem21_BID),
    .m00_axi_bready(m_axi_rmem21_BREADY),
    .m00_axi_bresp(m_axi_rmem21_BRESP),
    .m00_axi_bvalid(m_axi_rmem21_BVALID),
    .m00_axi_rdata(m_axi_rmem21_RDATA),
    .m00_axi_rid(m_axi_rmem21_RID),
    .m00_axi_rlast(m_axi_rmem21_RLAST),
    .m00_axi_rready(m_axi_rmem21_RREADY),
    .m00_axi_rresp(m_axi_rmem21_RRESP),
    .m00_axi_rvalid(m_axi_rmem21_RVALID),
    .m00_axi_wdata(m_axi_rmem21_WDATA),
    .m00_axi_wlast(m_axi_rmem21_WLAST),
    .m00_axi_wready(m_axi_rmem21_WREADY),
    .m00_axi_wstrb(m_axi_rmem21_WSTRB),
    .m00_axi_wvalid(m_axi_rmem21_WVALID),
    .s00_axi_araddr(m_axi_rmem21___Mmap2Stream_21___mmap_ARADDR),
    .s00_axi_arburst(m_axi_rmem21___Mmap2Stream_21___mmap_ARBURST),
    .s00_axi_arcache(m_axi_rmem21___Mmap2Stream_21___mmap_ARCACHE),
    .s00_axi_arid(m_axi_rmem21___Mmap2Stream_21___mmap_ARID),
    .s00_axi_arlen(m_axi_rmem21___Mmap2Stream_21___mmap_ARLEN),
    .s00_axi_arlock(m_axi_rmem21___Mmap2Stream_21___mmap_ARLOCK),
    .s00_axi_arprot(m_axi_rmem21___Mmap2Stream_21___mmap_ARPROT),
    .s00_axi_arqos(m_axi_rmem21___Mmap2Stream_21___mmap_ARQOS),
    .s00_axi_arready(m_axi_rmem21___Mmap2Stream_21___mmap_ARREADY),
    .s00_axi_arsize(m_axi_rmem21___Mmap2Stream_21___mmap_ARSIZE),
    .s00_axi_arvalid(m_axi_rmem21___Mmap2Stream_21___mmap_ARVALID),
    .s00_axi_awaddr(m_axi_rmem21___Mmap2Stream_21___mmap_AWADDR),
    .s00_axi_awburst(m_axi_rmem21___Mmap2Stream_21___mmap_AWBURST),
    .s00_axi_awcache(m_axi_rmem21___Mmap2Stream_21___mmap_AWCACHE),
    .s00_axi_awid(m_axi_rmem21___Mmap2Stream_21___mmap_AWID),
    .s00_axi_awlen(m_axi_rmem21___Mmap2Stream_21___mmap_AWLEN),
    .s00_axi_awlock(m_axi_rmem21___Mmap2Stream_21___mmap_AWLOCK),
    .s00_axi_awprot(m_axi_rmem21___Mmap2Stream_21___mmap_AWPROT),
    .s00_axi_awqos(m_axi_rmem21___Mmap2Stream_21___mmap_AWQOS),
    .s00_axi_awready(m_axi_rmem21___Mmap2Stream_21___mmap_AWREADY),
    .s00_axi_awsize(m_axi_rmem21___Mmap2Stream_21___mmap_AWSIZE),
    .s00_axi_awvalid(m_axi_rmem21___Mmap2Stream_21___mmap_AWVALID),
    .s00_axi_bid(m_axi_rmem21___Mmap2Stream_21___mmap_BID),
    .s00_axi_bready(m_axi_rmem21___Mmap2Stream_21___mmap_BREADY),
    .s00_axi_bresp(m_axi_rmem21___Mmap2Stream_21___mmap_BRESP),
    .s00_axi_bvalid(m_axi_rmem21___Mmap2Stream_21___mmap_BVALID),
    .s00_axi_rdata(m_axi_rmem21___Mmap2Stream_21___mmap_RDATA),
    .s00_axi_rid(m_axi_rmem21___Mmap2Stream_21___mmap_RID),
    .s00_axi_rlast(m_axi_rmem21___Mmap2Stream_21___mmap_RLAST),
    .s00_axi_rready(m_axi_rmem21___Mmap2Stream_21___mmap_RREADY),
    .s00_axi_rresp(m_axi_rmem21___Mmap2Stream_21___mmap_RRESP),
    .s00_axi_rvalid(m_axi_rmem21___Mmap2Stream_21___mmap_RVALID),
    .s00_axi_wdata(m_axi_rmem21___Mmap2Stream_21___mmap_WDATA),
    .s00_axi_wlast(m_axi_rmem21___Mmap2Stream_21___mmap_WLAST),
    .s00_axi_wready(m_axi_rmem21___Mmap2Stream_21___mmap_WREADY),
    .s00_axi_wstrb(m_axi_rmem21___Mmap2Stream_21___mmap_WSTRB),
    .s00_axi_wvalid(m_axi_rmem21___Mmap2Stream_21___mmap_WVALID),
    .s01_axi_araddr(m_axi_rmem21___Stream2Mmap_21___mmap_ARADDR),
    .s01_axi_arburst(m_axi_rmem21___Stream2Mmap_21___mmap_ARBURST),
    .s01_axi_arcache(m_axi_rmem21___Stream2Mmap_21___mmap_ARCACHE),
    .s01_axi_arid(m_axi_rmem21___Stream2Mmap_21___mmap_ARID),
    .s01_axi_arlen(m_axi_rmem21___Stream2Mmap_21___mmap_ARLEN),
    .s01_axi_arlock(m_axi_rmem21___Stream2Mmap_21___mmap_ARLOCK),
    .s01_axi_arprot(m_axi_rmem21___Stream2Mmap_21___mmap_ARPROT),
    .s01_axi_arqos(m_axi_rmem21___Stream2Mmap_21___mmap_ARQOS),
    .s01_axi_arready(m_axi_rmem21___Stream2Mmap_21___mmap_ARREADY),
    .s01_axi_arsize(m_axi_rmem21___Stream2Mmap_21___mmap_ARSIZE),
    .s01_axi_arvalid(m_axi_rmem21___Stream2Mmap_21___mmap_ARVALID),
    .s01_axi_awaddr(m_axi_rmem21___Stream2Mmap_21___mmap_AWADDR),
    .s01_axi_awburst(m_axi_rmem21___Stream2Mmap_21___mmap_AWBURST),
    .s01_axi_awcache(m_axi_rmem21___Stream2Mmap_21___mmap_AWCACHE),
    .s01_axi_awid(m_axi_rmem21___Stream2Mmap_21___mmap_AWID),
    .s01_axi_awlen(m_axi_rmem21___Stream2Mmap_21___mmap_AWLEN),
    .s01_axi_awlock(m_axi_rmem21___Stream2Mmap_21___mmap_AWLOCK),
    .s01_axi_awprot(m_axi_rmem21___Stream2Mmap_21___mmap_AWPROT),
    .s01_axi_awqos(m_axi_rmem21___Stream2Mmap_21___mmap_AWQOS),
    .s01_axi_awready(m_axi_rmem21___Stream2Mmap_21___mmap_AWREADY),
    .s01_axi_awsize(m_axi_rmem21___Stream2Mmap_21___mmap_AWSIZE),
    .s01_axi_awvalid(m_axi_rmem21___Stream2Mmap_21___mmap_AWVALID),
    .s01_axi_bid(m_axi_rmem21___Stream2Mmap_21___mmap_BID),
    .s01_axi_bready(m_axi_rmem21___Stream2Mmap_21___mmap_BREADY),
    .s01_axi_bresp(m_axi_rmem21___Stream2Mmap_21___mmap_BRESP),
    .s01_axi_bvalid(m_axi_rmem21___Stream2Mmap_21___mmap_BVALID),
    .s01_axi_rdata(m_axi_rmem21___Stream2Mmap_21___mmap_RDATA),
    .s01_axi_rid(m_axi_rmem21___Stream2Mmap_21___mmap_RID),
    .s01_axi_rlast(m_axi_rmem21___Stream2Mmap_21___mmap_RLAST),
    .s01_axi_rready(m_axi_rmem21___Stream2Mmap_21___mmap_RREADY),
    .s01_axi_rresp(m_axi_rmem21___Stream2Mmap_21___mmap_RRESP),
    .s01_axi_rvalid(m_axi_rmem21___Stream2Mmap_21___mmap_RVALID),
    .s01_axi_wdata(m_axi_rmem21___Stream2Mmap_21___mmap_WDATA),
    .s01_axi_wlast(m_axi_rmem21___Stream2Mmap_21___mmap_WLAST),
    .s01_axi_wready(m_axi_rmem21___Stream2Mmap_21___mmap_WREADY),
    .s01_axi_wstrb(m_axi_rmem21___Stream2Mmap_21___mmap_WSTRB),
    .s01_axi_wvalid(m_axi_rmem21___Stream2Mmap_21___mmap_WVALID)
  );


  (* keep_hierarchy = "yes" *) axi_crossbar_2x1
  #(
    .DATA_WIDTH(512),
    .ADDR_WIDTH(64),
    .S_ID_WIDTH(1),
    .M_ID_WIDTH(2),
    .M00_ADDR_WIDTH(64),
    .M00_ISSUE(16),
    .S00_THREADS(1),
    .S01_THREADS(1)
  )
  axi_crossbar_2x1__rmem22
  (
    .clk(ap_clk),
    .rst(ap_rst_n_inv),
    .m00_axi_araddr(m_axi_rmem22_ARADDR),
    .m00_axi_arburst(m_axi_rmem22_ARBURST),
    .m00_axi_arcache(m_axi_rmem22_ARCACHE),
    .m00_axi_arid(m_axi_rmem22_ARID),
    .m00_axi_arlen(m_axi_rmem22_ARLEN),
    .m00_axi_arlock(m_axi_rmem22_ARLOCK),
    .m00_axi_arprot(m_axi_rmem22_ARPROT),
    .m00_axi_arqos(m_axi_rmem22_ARQOS),
    .m00_axi_arready(m_axi_rmem22_ARREADY),
    .m00_axi_arsize(m_axi_rmem22_ARSIZE),
    .m00_axi_arvalid(m_axi_rmem22_ARVALID),
    .m00_axi_awaddr(m_axi_rmem22_AWADDR),
    .m00_axi_awburst(m_axi_rmem22_AWBURST),
    .m00_axi_awcache(m_axi_rmem22_AWCACHE),
    .m00_axi_awid(m_axi_rmem22_AWID),
    .m00_axi_awlen(m_axi_rmem22_AWLEN),
    .m00_axi_awlock(m_axi_rmem22_AWLOCK),
    .m00_axi_awprot(m_axi_rmem22_AWPROT),
    .m00_axi_awqos(m_axi_rmem22_AWQOS),
    .m00_axi_awready(m_axi_rmem22_AWREADY),
    .m00_axi_awsize(m_axi_rmem22_AWSIZE),
    .m00_axi_awvalid(m_axi_rmem22_AWVALID),
    .m00_axi_bid(m_axi_rmem22_BID),
    .m00_axi_bready(m_axi_rmem22_BREADY),
    .m00_axi_bresp(m_axi_rmem22_BRESP),
    .m00_axi_bvalid(m_axi_rmem22_BVALID),
    .m00_axi_rdata(m_axi_rmem22_RDATA),
    .m00_axi_rid(m_axi_rmem22_RID),
    .m00_axi_rlast(m_axi_rmem22_RLAST),
    .m00_axi_rready(m_axi_rmem22_RREADY),
    .m00_axi_rresp(m_axi_rmem22_RRESP),
    .m00_axi_rvalid(m_axi_rmem22_RVALID),
    .m00_axi_wdata(m_axi_rmem22_WDATA),
    .m00_axi_wlast(m_axi_rmem22_WLAST),
    .m00_axi_wready(m_axi_rmem22_WREADY),
    .m00_axi_wstrb(m_axi_rmem22_WSTRB),
    .m00_axi_wvalid(m_axi_rmem22_WVALID),
    .s00_axi_araddr(m_axi_rmem22___Mmap2Stream_22___mmap_ARADDR),
    .s00_axi_arburst(m_axi_rmem22___Mmap2Stream_22___mmap_ARBURST),
    .s00_axi_arcache(m_axi_rmem22___Mmap2Stream_22___mmap_ARCACHE),
    .s00_axi_arid(m_axi_rmem22___Mmap2Stream_22___mmap_ARID),
    .s00_axi_arlen(m_axi_rmem22___Mmap2Stream_22___mmap_ARLEN),
    .s00_axi_arlock(m_axi_rmem22___Mmap2Stream_22___mmap_ARLOCK),
    .s00_axi_arprot(m_axi_rmem22___Mmap2Stream_22___mmap_ARPROT),
    .s00_axi_arqos(m_axi_rmem22___Mmap2Stream_22___mmap_ARQOS),
    .s00_axi_arready(m_axi_rmem22___Mmap2Stream_22___mmap_ARREADY),
    .s00_axi_arsize(m_axi_rmem22___Mmap2Stream_22___mmap_ARSIZE),
    .s00_axi_arvalid(m_axi_rmem22___Mmap2Stream_22___mmap_ARVALID),
    .s00_axi_awaddr(m_axi_rmem22___Mmap2Stream_22___mmap_AWADDR),
    .s00_axi_awburst(m_axi_rmem22___Mmap2Stream_22___mmap_AWBURST),
    .s00_axi_awcache(m_axi_rmem22___Mmap2Stream_22___mmap_AWCACHE),
    .s00_axi_awid(m_axi_rmem22___Mmap2Stream_22___mmap_AWID),
    .s00_axi_awlen(m_axi_rmem22___Mmap2Stream_22___mmap_AWLEN),
    .s00_axi_awlock(m_axi_rmem22___Mmap2Stream_22___mmap_AWLOCK),
    .s00_axi_awprot(m_axi_rmem22___Mmap2Stream_22___mmap_AWPROT),
    .s00_axi_awqos(m_axi_rmem22___Mmap2Stream_22___mmap_AWQOS),
    .s00_axi_awready(m_axi_rmem22___Mmap2Stream_22___mmap_AWREADY),
    .s00_axi_awsize(m_axi_rmem22___Mmap2Stream_22___mmap_AWSIZE),
    .s00_axi_awvalid(m_axi_rmem22___Mmap2Stream_22___mmap_AWVALID),
    .s00_axi_bid(m_axi_rmem22___Mmap2Stream_22___mmap_BID),
    .s00_axi_bready(m_axi_rmem22___Mmap2Stream_22___mmap_BREADY),
    .s00_axi_bresp(m_axi_rmem22___Mmap2Stream_22___mmap_BRESP),
    .s00_axi_bvalid(m_axi_rmem22___Mmap2Stream_22___mmap_BVALID),
    .s00_axi_rdata(m_axi_rmem22___Mmap2Stream_22___mmap_RDATA),
    .s00_axi_rid(m_axi_rmem22___Mmap2Stream_22___mmap_RID),
    .s00_axi_rlast(m_axi_rmem22___Mmap2Stream_22___mmap_RLAST),
    .s00_axi_rready(m_axi_rmem22___Mmap2Stream_22___mmap_RREADY),
    .s00_axi_rresp(m_axi_rmem22___Mmap2Stream_22___mmap_RRESP),
    .s00_axi_rvalid(m_axi_rmem22___Mmap2Stream_22___mmap_RVALID),
    .s00_axi_wdata(m_axi_rmem22___Mmap2Stream_22___mmap_WDATA),
    .s00_axi_wlast(m_axi_rmem22___Mmap2Stream_22___mmap_WLAST),
    .s00_axi_wready(m_axi_rmem22___Mmap2Stream_22___mmap_WREADY),
    .s00_axi_wstrb(m_axi_rmem22___Mmap2Stream_22___mmap_WSTRB),
    .s00_axi_wvalid(m_axi_rmem22___Mmap2Stream_22___mmap_WVALID),
    .s01_axi_araddr(m_axi_rmem22___Stream2Mmap_22___mmap_ARADDR),
    .s01_axi_arburst(m_axi_rmem22___Stream2Mmap_22___mmap_ARBURST),
    .s01_axi_arcache(m_axi_rmem22___Stream2Mmap_22___mmap_ARCACHE),
    .s01_axi_arid(m_axi_rmem22___Stream2Mmap_22___mmap_ARID),
    .s01_axi_arlen(m_axi_rmem22___Stream2Mmap_22___mmap_ARLEN),
    .s01_axi_arlock(m_axi_rmem22___Stream2Mmap_22___mmap_ARLOCK),
    .s01_axi_arprot(m_axi_rmem22___Stream2Mmap_22___mmap_ARPROT),
    .s01_axi_arqos(m_axi_rmem22___Stream2Mmap_22___mmap_ARQOS),
    .s01_axi_arready(m_axi_rmem22___Stream2Mmap_22___mmap_ARREADY),
    .s01_axi_arsize(m_axi_rmem22___Stream2Mmap_22___mmap_ARSIZE),
    .s01_axi_arvalid(m_axi_rmem22___Stream2Mmap_22___mmap_ARVALID),
    .s01_axi_awaddr(m_axi_rmem22___Stream2Mmap_22___mmap_AWADDR),
    .s01_axi_awburst(m_axi_rmem22___Stream2Mmap_22___mmap_AWBURST),
    .s01_axi_awcache(m_axi_rmem22___Stream2Mmap_22___mmap_AWCACHE),
    .s01_axi_awid(m_axi_rmem22___Stream2Mmap_22___mmap_AWID),
    .s01_axi_awlen(m_axi_rmem22___Stream2Mmap_22___mmap_AWLEN),
    .s01_axi_awlock(m_axi_rmem22___Stream2Mmap_22___mmap_AWLOCK),
    .s01_axi_awprot(m_axi_rmem22___Stream2Mmap_22___mmap_AWPROT),
    .s01_axi_awqos(m_axi_rmem22___Stream2Mmap_22___mmap_AWQOS),
    .s01_axi_awready(m_axi_rmem22___Stream2Mmap_22___mmap_AWREADY),
    .s01_axi_awsize(m_axi_rmem22___Stream2Mmap_22___mmap_AWSIZE),
    .s01_axi_awvalid(m_axi_rmem22___Stream2Mmap_22___mmap_AWVALID),
    .s01_axi_bid(m_axi_rmem22___Stream2Mmap_22___mmap_BID),
    .s01_axi_bready(m_axi_rmem22___Stream2Mmap_22___mmap_BREADY),
    .s01_axi_bresp(m_axi_rmem22___Stream2Mmap_22___mmap_BRESP),
    .s01_axi_bvalid(m_axi_rmem22___Stream2Mmap_22___mmap_BVALID),
    .s01_axi_rdata(m_axi_rmem22___Stream2Mmap_22___mmap_RDATA),
    .s01_axi_rid(m_axi_rmem22___Stream2Mmap_22___mmap_RID),
    .s01_axi_rlast(m_axi_rmem22___Stream2Mmap_22___mmap_RLAST),
    .s01_axi_rready(m_axi_rmem22___Stream2Mmap_22___mmap_RREADY),
    .s01_axi_rresp(m_axi_rmem22___Stream2Mmap_22___mmap_RRESP),
    .s01_axi_rvalid(m_axi_rmem22___Stream2Mmap_22___mmap_RVALID),
    .s01_axi_wdata(m_axi_rmem22___Stream2Mmap_22___mmap_WDATA),
    .s01_axi_wlast(m_axi_rmem22___Stream2Mmap_22___mmap_WLAST),
    .s01_axi_wready(m_axi_rmem22___Stream2Mmap_22___mmap_WREADY),
    .s01_axi_wstrb(m_axi_rmem22___Stream2Mmap_22___mmap_WSTRB),
    .s01_axi_wvalid(m_axi_rmem22___Stream2Mmap_22___mmap_WVALID)
  );


  (* keep_hierarchy = "yes" *) axi_crossbar_2x1
  #(
    .DATA_WIDTH(512),
    .ADDR_WIDTH(64),
    .S_ID_WIDTH(1),
    .M_ID_WIDTH(2),
    .M00_ADDR_WIDTH(64),
    .M00_ISSUE(16),
    .S00_THREADS(1),
    .S01_THREADS(1)
  )
  axi_crossbar_2x1__rmem23
  (
    .clk(ap_clk),
    .rst(ap_rst_n_inv),
    .m00_axi_araddr(m_axi_rmem23_ARADDR),
    .m00_axi_arburst(m_axi_rmem23_ARBURST),
    .m00_axi_arcache(m_axi_rmem23_ARCACHE),
    .m00_axi_arid(m_axi_rmem23_ARID),
    .m00_axi_arlen(m_axi_rmem23_ARLEN),
    .m00_axi_arlock(m_axi_rmem23_ARLOCK),
    .m00_axi_arprot(m_axi_rmem23_ARPROT),
    .m00_axi_arqos(m_axi_rmem23_ARQOS),
    .m00_axi_arready(m_axi_rmem23_ARREADY),
    .m00_axi_arsize(m_axi_rmem23_ARSIZE),
    .m00_axi_arvalid(m_axi_rmem23_ARVALID),
    .m00_axi_awaddr(m_axi_rmem23_AWADDR),
    .m00_axi_awburst(m_axi_rmem23_AWBURST),
    .m00_axi_awcache(m_axi_rmem23_AWCACHE),
    .m00_axi_awid(m_axi_rmem23_AWID),
    .m00_axi_awlen(m_axi_rmem23_AWLEN),
    .m00_axi_awlock(m_axi_rmem23_AWLOCK),
    .m00_axi_awprot(m_axi_rmem23_AWPROT),
    .m00_axi_awqos(m_axi_rmem23_AWQOS),
    .m00_axi_awready(m_axi_rmem23_AWREADY),
    .m00_axi_awsize(m_axi_rmem23_AWSIZE),
    .m00_axi_awvalid(m_axi_rmem23_AWVALID),
    .m00_axi_bid(m_axi_rmem23_BID),
    .m00_axi_bready(m_axi_rmem23_BREADY),
    .m00_axi_bresp(m_axi_rmem23_BRESP),
    .m00_axi_bvalid(m_axi_rmem23_BVALID),
    .m00_axi_rdata(m_axi_rmem23_RDATA),
    .m00_axi_rid(m_axi_rmem23_RID),
    .m00_axi_rlast(m_axi_rmem23_RLAST),
    .m00_axi_rready(m_axi_rmem23_RREADY),
    .m00_axi_rresp(m_axi_rmem23_RRESP),
    .m00_axi_rvalid(m_axi_rmem23_RVALID),
    .m00_axi_wdata(m_axi_rmem23_WDATA),
    .m00_axi_wlast(m_axi_rmem23_WLAST),
    .m00_axi_wready(m_axi_rmem23_WREADY),
    .m00_axi_wstrb(m_axi_rmem23_WSTRB),
    .m00_axi_wvalid(m_axi_rmem23_WVALID),
    .s00_axi_araddr(m_axi_rmem23___Mmap2Stream_23___mmap_ARADDR),
    .s00_axi_arburst(m_axi_rmem23___Mmap2Stream_23___mmap_ARBURST),
    .s00_axi_arcache(m_axi_rmem23___Mmap2Stream_23___mmap_ARCACHE),
    .s00_axi_arid(m_axi_rmem23___Mmap2Stream_23___mmap_ARID),
    .s00_axi_arlen(m_axi_rmem23___Mmap2Stream_23___mmap_ARLEN),
    .s00_axi_arlock(m_axi_rmem23___Mmap2Stream_23___mmap_ARLOCK),
    .s00_axi_arprot(m_axi_rmem23___Mmap2Stream_23___mmap_ARPROT),
    .s00_axi_arqos(m_axi_rmem23___Mmap2Stream_23___mmap_ARQOS),
    .s00_axi_arready(m_axi_rmem23___Mmap2Stream_23___mmap_ARREADY),
    .s00_axi_arsize(m_axi_rmem23___Mmap2Stream_23___mmap_ARSIZE),
    .s00_axi_arvalid(m_axi_rmem23___Mmap2Stream_23___mmap_ARVALID),
    .s00_axi_awaddr(m_axi_rmem23___Mmap2Stream_23___mmap_AWADDR),
    .s00_axi_awburst(m_axi_rmem23___Mmap2Stream_23___mmap_AWBURST),
    .s00_axi_awcache(m_axi_rmem23___Mmap2Stream_23___mmap_AWCACHE),
    .s00_axi_awid(m_axi_rmem23___Mmap2Stream_23___mmap_AWID),
    .s00_axi_awlen(m_axi_rmem23___Mmap2Stream_23___mmap_AWLEN),
    .s00_axi_awlock(m_axi_rmem23___Mmap2Stream_23___mmap_AWLOCK),
    .s00_axi_awprot(m_axi_rmem23___Mmap2Stream_23___mmap_AWPROT),
    .s00_axi_awqos(m_axi_rmem23___Mmap2Stream_23___mmap_AWQOS),
    .s00_axi_awready(m_axi_rmem23___Mmap2Stream_23___mmap_AWREADY),
    .s00_axi_awsize(m_axi_rmem23___Mmap2Stream_23___mmap_AWSIZE),
    .s00_axi_awvalid(m_axi_rmem23___Mmap2Stream_23___mmap_AWVALID),
    .s00_axi_bid(m_axi_rmem23___Mmap2Stream_23___mmap_BID),
    .s00_axi_bready(m_axi_rmem23___Mmap2Stream_23___mmap_BREADY),
    .s00_axi_bresp(m_axi_rmem23___Mmap2Stream_23___mmap_BRESP),
    .s00_axi_bvalid(m_axi_rmem23___Mmap2Stream_23___mmap_BVALID),
    .s00_axi_rdata(m_axi_rmem23___Mmap2Stream_23___mmap_RDATA),
    .s00_axi_rid(m_axi_rmem23___Mmap2Stream_23___mmap_RID),
    .s00_axi_rlast(m_axi_rmem23___Mmap2Stream_23___mmap_RLAST),
    .s00_axi_rready(m_axi_rmem23___Mmap2Stream_23___mmap_RREADY),
    .s00_axi_rresp(m_axi_rmem23___Mmap2Stream_23___mmap_RRESP),
    .s00_axi_rvalid(m_axi_rmem23___Mmap2Stream_23___mmap_RVALID),
    .s00_axi_wdata(m_axi_rmem23___Mmap2Stream_23___mmap_WDATA),
    .s00_axi_wlast(m_axi_rmem23___Mmap2Stream_23___mmap_WLAST),
    .s00_axi_wready(m_axi_rmem23___Mmap2Stream_23___mmap_WREADY),
    .s00_axi_wstrb(m_axi_rmem23___Mmap2Stream_23___mmap_WSTRB),
    .s00_axi_wvalid(m_axi_rmem23___Mmap2Stream_23___mmap_WVALID),
    .s01_axi_araddr(m_axi_rmem23___Stream2Mmap_23___mmap_ARADDR),
    .s01_axi_arburst(m_axi_rmem23___Stream2Mmap_23___mmap_ARBURST),
    .s01_axi_arcache(m_axi_rmem23___Stream2Mmap_23___mmap_ARCACHE),
    .s01_axi_arid(m_axi_rmem23___Stream2Mmap_23___mmap_ARID),
    .s01_axi_arlen(m_axi_rmem23___Stream2Mmap_23___mmap_ARLEN),
    .s01_axi_arlock(m_axi_rmem23___Stream2Mmap_23___mmap_ARLOCK),
    .s01_axi_arprot(m_axi_rmem23___Stream2Mmap_23___mmap_ARPROT),
    .s01_axi_arqos(m_axi_rmem23___Stream2Mmap_23___mmap_ARQOS),
    .s01_axi_arready(m_axi_rmem23___Stream2Mmap_23___mmap_ARREADY),
    .s01_axi_arsize(m_axi_rmem23___Stream2Mmap_23___mmap_ARSIZE),
    .s01_axi_arvalid(m_axi_rmem23___Stream2Mmap_23___mmap_ARVALID),
    .s01_axi_awaddr(m_axi_rmem23___Stream2Mmap_23___mmap_AWADDR),
    .s01_axi_awburst(m_axi_rmem23___Stream2Mmap_23___mmap_AWBURST),
    .s01_axi_awcache(m_axi_rmem23___Stream2Mmap_23___mmap_AWCACHE),
    .s01_axi_awid(m_axi_rmem23___Stream2Mmap_23___mmap_AWID),
    .s01_axi_awlen(m_axi_rmem23___Stream2Mmap_23___mmap_AWLEN),
    .s01_axi_awlock(m_axi_rmem23___Stream2Mmap_23___mmap_AWLOCK),
    .s01_axi_awprot(m_axi_rmem23___Stream2Mmap_23___mmap_AWPROT),
    .s01_axi_awqos(m_axi_rmem23___Stream2Mmap_23___mmap_AWQOS),
    .s01_axi_awready(m_axi_rmem23___Stream2Mmap_23___mmap_AWREADY),
    .s01_axi_awsize(m_axi_rmem23___Stream2Mmap_23___mmap_AWSIZE),
    .s01_axi_awvalid(m_axi_rmem23___Stream2Mmap_23___mmap_AWVALID),
    .s01_axi_bid(m_axi_rmem23___Stream2Mmap_23___mmap_BID),
    .s01_axi_bready(m_axi_rmem23___Stream2Mmap_23___mmap_BREADY),
    .s01_axi_bresp(m_axi_rmem23___Stream2Mmap_23___mmap_BRESP),
    .s01_axi_bvalid(m_axi_rmem23___Stream2Mmap_23___mmap_BVALID),
    .s01_axi_rdata(m_axi_rmem23___Stream2Mmap_23___mmap_RDATA),
    .s01_axi_rid(m_axi_rmem23___Stream2Mmap_23___mmap_RID),
    .s01_axi_rlast(m_axi_rmem23___Stream2Mmap_23___mmap_RLAST),
    .s01_axi_rready(m_axi_rmem23___Stream2Mmap_23___mmap_RREADY),
    .s01_axi_rresp(m_axi_rmem23___Stream2Mmap_23___mmap_RRESP),
    .s01_axi_rvalid(m_axi_rmem23___Stream2Mmap_23___mmap_RVALID),
    .s01_axi_wdata(m_axi_rmem23___Stream2Mmap_23___mmap_WDATA),
    .s01_axi_wlast(m_axi_rmem23___Stream2Mmap_23___mmap_WLAST),
    .s01_axi_wready(m_axi_rmem23___Stream2Mmap_23___mmap_WREADY),
    .s01_axi_wstrb(m_axi_rmem23___Stream2Mmap_23___mmap_WSTRB),
    .s01_axi_wvalid(m_axi_rmem23___Stream2Mmap_23___mmap_WVALID)
  );


  (* keep_hierarchy = "yes" *) axi_crossbar_2x1
  #(
    .DATA_WIDTH(512),
    .ADDR_WIDTH(64),
    .S_ID_WIDTH(1),
    .M_ID_WIDTH(2),
    .M00_ADDR_WIDTH(64),
    .M00_ISSUE(16),
    .S00_THREADS(1),
    .S01_THREADS(1)
  )
  axi_crossbar_2x1__rmem24
  (
    .clk(ap_clk),
    .rst(ap_rst_n_inv),
    .m00_axi_araddr(m_axi_rmem24_ARADDR),
    .m00_axi_arburst(m_axi_rmem24_ARBURST),
    .m00_axi_arcache(m_axi_rmem24_ARCACHE),
    .m00_axi_arid(m_axi_rmem24_ARID),
    .m00_axi_arlen(m_axi_rmem24_ARLEN),
    .m00_axi_arlock(m_axi_rmem24_ARLOCK),
    .m00_axi_arprot(m_axi_rmem24_ARPROT),
    .m00_axi_arqos(m_axi_rmem24_ARQOS),
    .m00_axi_arready(m_axi_rmem24_ARREADY),
    .m00_axi_arsize(m_axi_rmem24_ARSIZE),
    .m00_axi_arvalid(m_axi_rmem24_ARVALID),
    .m00_axi_awaddr(m_axi_rmem24_AWADDR),
    .m00_axi_awburst(m_axi_rmem24_AWBURST),
    .m00_axi_awcache(m_axi_rmem24_AWCACHE),
    .m00_axi_awid(m_axi_rmem24_AWID),
    .m00_axi_awlen(m_axi_rmem24_AWLEN),
    .m00_axi_awlock(m_axi_rmem24_AWLOCK),
    .m00_axi_awprot(m_axi_rmem24_AWPROT),
    .m00_axi_awqos(m_axi_rmem24_AWQOS),
    .m00_axi_awready(m_axi_rmem24_AWREADY),
    .m00_axi_awsize(m_axi_rmem24_AWSIZE),
    .m00_axi_awvalid(m_axi_rmem24_AWVALID),
    .m00_axi_bid(m_axi_rmem24_BID),
    .m00_axi_bready(m_axi_rmem24_BREADY),
    .m00_axi_bresp(m_axi_rmem24_BRESP),
    .m00_axi_bvalid(m_axi_rmem24_BVALID),
    .m00_axi_rdata(m_axi_rmem24_RDATA),
    .m00_axi_rid(m_axi_rmem24_RID),
    .m00_axi_rlast(m_axi_rmem24_RLAST),
    .m00_axi_rready(m_axi_rmem24_RREADY),
    .m00_axi_rresp(m_axi_rmem24_RRESP),
    .m00_axi_rvalid(m_axi_rmem24_RVALID),
    .m00_axi_wdata(m_axi_rmem24_WDATA),
    .m00_axi_wlast(m_axi_rmem24_WLAST),
    .m00_axi_wready(m_axi_rmem24_WREADY),
    .m00_axi_wstrb(m_axi_rmem24_WSTRB),
    .m00_axi_wvalid(m_axi_rmem24_WVALID),
    .s00_axi_araddr(m_axi_rmem24___Mmap2Stream_24___mmap_ARADDR),
    .s00_axi_arburst(m_axi_rmem24___Mmap2Stream_24___mmap_ARBURST),
    .s00_axi_arcache(m_axi_rmem24___Mmap2Stream_24___mmap_ARCACHE),
    .s00_axi_arid(m_axi_rmem24___Mmap2Stream_24___mmap_ARID),
    .s00_axi_arlen(m_axi_rmem24___Mmap2Stream_24___mmap_ARLEN),
    .s00_axi_arlock(m_axi_rmem24___Mmap2Stream_24___mmap_ARLOCK),
    .s00_axi_arprot(m_axi_rmem24___Mmap2Stream_24___mmap_ARPROT),
    .s00_axi_arqos(m_axi_rmem24___Mmap2Stream_24___mmap_ARQOS),
    .s00_axi_arready(m_axi_rmem24___Mmap2Stream_24___mmap_ARREADY),
    .s00_axi_arsize(m_axi_rmem24___Mmap2Stream_24___mmap_ARSIZE),
    .s00_axi_arvalid(m_axi_rmem24___Mmap2Stream_24___mmap_ARVALID),
    .s00_axi_awaddr(m_axi_rmem24___Mmap2Stream_24___mmap_AWADDR),
    .s00_axi_awburst(m_axi_rmem24___Mmap2Stream_24___mmap_AWBURST),
    .s00_axi_awcache(m_axi_rmem24___Mmap2Stream_24___mmap_AWCACHE),
    .s00_axi_awid(m_axi_rmem24___Mmap2Stream_24___mmap_AWID),
    .s00_axi_awlen(m_axi_rmem24___Mmap2Stream_24___mmap_AWLEN),
    .s00_axi_awlock(m_axi_rmem24___Mmap2Stream_24___mmap_AWLOCK),
    .s00_axi_awprot(m_axi_rmem24___Mmap2Stream_24___mmap_AWPROT),
    .s00_axi_awqos(m_axi_rmem24___Mmap2Stream_24___mmap_AWQOS),
    .s00_axi_awready(m_axi_rmem24___Mmap2Stream_24___mmap_AWREADY),
    .s00_axi_awsize(m_axi_rmem24___Mmap2Stream_24___mmap_AWSIZE),
    .s00_axi_awvalid(m_axi_rmem24___Mmap2Stream_24___mmap_AWVALID),
    .s00_axi_bid(m_axi_rmem24___Mmap2Stream_24___mmap_BID),
    .s00_axi_bready(m_axi_rmem24___Mmap2Stream_24___mmap_BREADY),
    .s00_axi_bresp(m_axi_rmem24___Mmap2Stream_24___mmap_BRESP),
    .s00_axi_bvalid(m_axi_rmem24___Mmap2Stream_24___mmap_BVALID),
    .s00_axi_rdata(m_axi_rmem24___Mmap2Stream_24___mmap_RDATA),
    .s00_axi_rid(m_axi_rmem24___Mmap2Stream_24___mmap_RID),
    .s00_axi_rlast(m_axi_rmem24___Mmap2Stream_24___mmap_RLAST),
    .s00_axi_rready(m_axi_rmem24___Mmap2Stream_24___mmap_RREADY),
    .s00_axi_rresp(m_axi_rmem24___Mmap2Stream_24___mmap_RRESP),
    .s00_axi_rvalid(m_axi_rmem24___Mmap2Stream_24___mmap_RVALID),
    .s00_axi_wdata(m_axi_rmem24___Mmap2Stream_24___mmap_WDATA),
    .s00_axi_wlast(m_axi_rmem24___Mmap2Stream_24___mmap_WLAST),
    .s00_axi_wready(m_axi_rmem24___Mmap2Stream_24___mmap_WREADY),
    .s00_axi_wstrb(m_axi_rmem24___Mmap2Stream_24___mmap_WSTRB),
    .s00_axi_wvalid(m_axi_rmem24___Mmap2Stream_24___mmap_WVALID),
    .s01_axi_araddr(m_axi_rmem24___Stream2Mmap_24___mmap_ARADDR),
    .s01_axi_arburst(m_axi_rmem24___Stream2Mmap_24___mmap_ARBURST),
    .s01_axi_arcache(m_axi_rmem24___Stream2Mmap_24___mmap_ARCACHE),
    .s01_axi_arid(m_axi_rmem24___Stream2Mmap_24___mmap_ARID),
    .s01_axi_arlen(m_axi_rmem24___Stream2Mmap_24___mmap_ARLEN),
    .s01_axi_arlock(m_axi_rmem24___Stream2Mmap_24___mmap_ARLOCK),
    .s01_axi_arprot(m_axi_rmem24___Stream2Mmap_24___mmap_ARPROT),
    .s01_axi_arqos(m_axi_rmem24___Stream2Mmap_24___mmap_ARQOS),
    .s01_axi_arready(m_axi_rmem24___Stream2Mmap_24___mmap_ARREADY),
    .s01_axi_arsize(m_axi_rmem24___Stream2Mmap_24___mmap_ARSIZE),
    .s01_axi_arvalid(m_axi_rmem24___Stream2Mmap_24___mmap_ARVALID),
    .s01_axi_awaddr(m_axi_rmem24___Stream2Mmap_24___mmap_AWADDR),
    .s01_axi_awburst(m_axi_rmem24___Stream2Mmap_24___mmap_AWBURST),
    .s01_axi_awcache(m_axi_rmem24___Stream2Mmap_24___mmap_AWCACHE),
    .s01_axi_awid(m_axi_rmem24___Stream2Mmap_24___mmap_AWID),
    .s01_axi_awlen(m_axi_rmem24___Stream2Mmap_24___mmap_AWLEN),
    .s01_axi_awlock(m_axi_rmem24___Stream2Mmap_24___mmap_AWLOCK),
    .s01_axi_awprot(m_axi_rmem24___Stream2Mmap_24___mmap_AWPROT),
    .s01_axi_awqos(m_axi_rmem24___Stream2Mmap_24___mmap_AWQOS),
    .s01_axi_awready(m_axi_rmem24___Stream2Mmap_24___mmap_AWREADY),
    .s01_axi_awsize(m_axi_rmem24___Stream2Mmap_24___mmap_AWSIZE),
    .s01_axi_awvalid(m_axi_rmem24___Stream2Mmap_24___mmap_AWVALID),
    .s01_axi_bid(m_axi_rmem24___Stream2Mmap_24___mmap_BID),
    .s01_axi_bready(m_axi_rmem24___Stream2Mmap_24___mmap_BREADY),
    .s01_axi_bresp(m_axi_rmem24___Stream2Mmap_24___mmap_BRESP),
    .s01_axi_bvalid(m_axi_rmem24___Stream2Mmap_24___mmap_BVALID),
    .s01_axi_rdata(m_axi_rmem24___Stream2Mmap_24___mmap_RDATA),
    .s01_axi_rid(m_axi_rmem24___Stream2Mmap_24___mmap_RID),
    .s01_axi_rlast(m_axi_rmem24___Stream2Mmap_24___mmap_RLAST),
    .s01_axi_rready(m_axi_rmem24___Stream2Mmap_24___mmap_RREADY),
    .s01_axi_rresp(m_axi_rmem24___Stream2Mmap_24___mmap_RRESP),
    .s01_axi_rvalid(m_axi_rmem24___Stream2Mmap_24___mmap_RVALID),
    .s01_axi_wdata(m_axi_rmem24___Stream2Mmap_24___mmap_WDATA),
    .s01_axi_wlast(m_axi_rmem24___Stream2Mmap_24___mmap_WLAST),
    .s01_axi_wready(m_axi_rmem24___Stream2Mmap_24___mmap_WREADY),
    .s01_axi_wstrb(m_axi_rmem24___Stream2Mmap_24___mmap_WSTRB),
    .s01_axi_wvalid(m_axi_rmem24___Stream2Mmap_24___mmap_WVALID)
  );


  (* keep_hierarchy = "yes" *) axi_crossbar_2x1
  #(
    .DATA_WIDTH(512),
    .ADDR_WIDTH(64),
    .S_ID_WIDTH(1),
    .M_ID_WIDTH(2),
    .M00_ADDR_WIDTH(64),
    .M00_ISSUE(16),
    .S00_THREADS(1),
    .S01_THREADS(1)
  )
  axi_crossbar_2x1__rmem25
  (
    .clk(ap_clk),
    .rst(ap_rst_n_inv),
    .m00_axi_araddr(m_axi_rmem25_ARADDR),
    .m00_axi_arburst(m_axi_rmem25_ARBURST),
    .m00_axi_arcache(m_axi_rmem25_ARCACHE),
    .m00_axi_arid(m_axi_rmem25_ARID),
    .m00_axi_arlen(m_axi_rmem25_ARLEN),
    .m00_axi_arlock(m_axi_rmem25_ARLOCK),
    .m00_axi_arprot(m_axi_rmem25_ARPROT),
    .m00_axi_arqos(m_axi_rmem25_ARQOS),
    .m00_axi_arready(m_axi_rmem25_ARREADY),
    .m00_axi_arsize(m_axi_rmem25_ARSIZE),
    .m00_axi_arvalid(m_axi_rmem25_ARVALID),
    .m00_axi_awaddr(m_axi_rmem25_AWADDR),
    .m00_axi_awburst(m_axi_rmem25_AWBURST),
    .m00_axi_awcache(m_axi_rmem25_AWCACHE),
    .m00_axi_awid(m_axi_rmem25_AWID),
    .m00_axi_awlen(m_axi_rmem25_AWLEN),
    .m00_axi_awlock(m_axi_rmem25_AWLOCK),
    .m00_axi_awprot(m_axi_rmem25_AWPROT),
    .m00_axi_awqos(m_axi_rmem25_AWQOS),
    .m00_axi_awready(m_axi_rmem25_AWREADY),
    .m00_axi_awsize(m_axi_rmem25_AWSIZE),
    .m00_axi_awvalid(m_axi_rmem25_AWVALID),
    .m00_axi_bid(m_axi_rmem25_BID),
    .m00_axi_bready(m_axi_rmem25_BREADY),
    .m00_axi_bresp(m_axi_rmem25_BRESP),
    .m00_axi_bvalid(m_axi_rmem25_BVALID),
    .m00_axi_rdata(m_axi_rmem25_RDATA),
    .m00_axi_rid(m_axi_rmem25_RID),
    .m00_axi_rlast(m_axi_rmem25_RLAST),
    .m00_axi_rready(m_axi_rmem25_RREADY),
    .m00_axi_rresp(m_axi_rmem25_RRESP),
    .m00_axi_rvalid(m_axi_rmem25_RVALID),
    .m00_axi_wdata(m_axi_rmem25_WDATA),
    .m00_axi_wlast(m_axi_rmem25_WLAST),
    .m00_axi_wready(m_axi_rmem25_WREADY),
    .m00_axi_wstrb(m_axi_rmem25_WSTRB),
    .m00_axi_wvalid(m_axi_rmem25_WVALID),
    .s00_axi_araddr(m_axi_rmem25___Mmap2Stream_25___mmap_ARADDR),
    .s00_axi_arburst(m_axi_rmem25___Mmap2Stream_25___mmap_ARBURST),
    .s00_axi_arcache(m_axi_rmem25___Mmap2Stream_25___mmap_ARCACHE),
    .s00_axi_arid(m_axi_rmem25___Mmap2Stream_25___mmap_ARID),
    .s00_axi_arlen(m_axi_rmem25___Mmap2Stream_25___mmap_ARLEN),
    .s00_axi_arlock(m_axi_rmem25___Mmap2Stream_25___mmap_ARLOCK),
    .s00_axi_arprot(m_axi_rmem25___Mmap2Stream_25___mmap_ARPROT),
    .s00_axi_arqos(m_axi_rmem25___Mmap2Stream_25___mmap_ARQOS),
    .s00_axi_arready(m_axi_rmem25___Mmap2Stream_25___mmap_ARREADY),
    .s00_axi_arsize(m_axi_rmem25___Mmap2Stream_25___mmap_ARSIZE),
    .s00_axi_arvalid(m_axi_rmem25___Mmap2Stream_25___mmap_ARVALID),
    .s00_axi_awaddr(m_axi_rmem25___Mmap2Stream_25___mmap_AWADDR),
    .s00_axi_awburst(m_axi_rmem25___Mmap2Stream_25___mmap_AWBURST),
    .s00_axi_awcache(m_axi_rmem25___Mmap2Stream_25___mmap_AWCACHE),
    .s00_axi_awid(m_axi_rmem25___Mmap2Stream_25___mmap_AWID),
    .s00_axi_awlen(m_axi_rmem25___Mmap2Stream_25___mmap_AWLEN),
    .s00_axi_awlock(m_axi_rmem25___Mmap2Stream_25___mmap_AWLOCK),
    .s00_axi_awprot(m_axi_rmem25___Mmap2Stream_25___mmap_AWPROT),
    .s00_axi_awqos(m_axi_rmem25___Mmap2Stream_25___mmap_AWQOS),
    .s00_axi_awready(m_axi_rmem25___Mmap2Stream_25___mmap_AWREADY),
    .s00_axi_awsize(m_axi_rmem25___Mmap2Stream_25___mmap_AWSIZE),
    .s00_axi_awvalid(m_axi_rmem25___Mmap2Stream_25___mmap_AWVALID),
    .s00_axi_bid(m_axi_rmem25___Mmap2Stream_25___mmap_BID),
    .s00_axi_bready(m_axi_rmem25___Mmap2Stream_25___mmap_BREADY),
    .s00_axi_bresp(m_axi_rmem25___Mmap2Stream_25___mmap_BRESP),
    .s00_axi_bvalid(m_axi_rmem25___Mmap2Stream_25___mmap_BVALID),
    .s00_axi_rdata(m_axi_rmem25___Mmap2Stream_25___mmap_RDATA),
    .s00_axi_rid(m_axi_rmem25___Mmap2Stream_25___mmap_RID),
    .s00_axi_rlast(m_axi_rmem25___Mmap2Stream_25___mmap_RLAST),
    .s00_axi_rready(m_axi_rmem25___Mmap2Stream_25___mmap_RREADY),
    .s00_axi_rresp(m_axi_rmem25___Mmap2Stream_25___mmap_RRESP),
    .s00_axi_rvalid(m_axi_rmem25___Mmap2Stream_25___mmap_RVALID),
    .s00_axi_wdata(m_axi_rmem25___Mmap2Stream_25___mmap_WDATA),
    .s00_axi_wlast(m_axi_rmem25___Mmap2Stream_25___mmap_WLAST),
    .s00_axi_wready(m_axi_rmem25___Mmap2Stream_25___mmap_WREADY),
    .s00_axi_wstrb(m_axi_rmem25___Mmap2Stream_25___mmap_WSTRB),
    .s00_axi_wvalid(m_axi_rmem25___Mmap2Stream_25___mmap_WVALID),
    .s01_axi_araddr(m_axi_rmem25___Stream2Mmap_25___mmap_ARADDR),
    .s01_axi_arburst(m_axi_rmem25___Stream2Mmap_25___mmap_ARBURST),
    .s01_axi_arcache(m_axi_rmem25___Stream2Mmap_25___mmap_ARCACHE),
    .s01_axi_arid(m_axi_rmem25___Stream2Mmap_25___mmap_ARID),
    .s01_axi_arlen(m_axi_rmem25___Stream2Mmap_25___mmap_ARLEN),
    .s01_axi_arlock(m_axi_rmem25___Stream2Mmap_25___mmap_ARLOCK),
    .s01_axi_arprot(m_axi_rmem25___Stream2Mmap_25___mmap_ARPROT),
    .s01_axi_arqos(m_axi_rmem25___Stream2Mmap_25___mmap_ARQOS),
    .s01_axi_arready(m_axi_rmem25___Stream2Mmap_25___mmap_ARREADY),
    .s01_axi_arsize(m_axi_rmem25___Stream2Mmap_25___mmap_ARSIZE),
    .s01_axi_arvalid(m_axi_rmem25___Stream2Mmap_25___mmap_ARVALID),
    .s01_axi_awaddr(m_axi_rmem25___Stream2Mmap_25___mmap_AWADDR),
    .s01_axi_awburst(m_axi_rmem25___Stream2Mmap_25___mmap_AWBURST),
    .s01_axi_awcache(m_axi_rmem25___Stream2Mmap_25___mmap_AWCACHE),
    .s01_axi_awid(m_axi_rmem25___Stream2Mmap_25___mmap_AWID),
    .s01_axi_awlen(m_axi_rmem25___Stream2Mmap_25___mmap_AWLEN),
    .s01_axi_awlock(m_axi_rmem25___Stream2Mmap_25___mmap_AWLOCK),
    .s01_axi_awprot(m_axi_rmem25___Stream2Mmap_25___mmap_AWPROT),
    .s01_axi_awqos(m_axi_rmem25___Stream2Mmap_25___mmap_AWQOS),
    .s01_axi_awready(m_axi_rmem25___Stream2Mmap_25___mmap_AWREADY),
    .s01_axi_awsize(m_axi_rmem25___Stream2Mmap_25___mmap_AWSIZE),
    .s01_axi_awvalid(m_axi_rmem25___Stream2Mmap_25___mmap_AWVALID),
    .s01_axi_bid(m_axi_rmem25___Stream2Mmap_25___mmap_BID),
    .s01_axi_bready(m_axi_rmem25___Stream2Mmap_25___mmap_BREADY),
    .s01_axi_bresp(m_axi_rmem25___Stream2Mmap_25___mmap_BRESP),
    .s01_axi_bvalid(m_axi_rmem25___Stream2Mmap_25___mmap_BVALID),
    .s01_axi_rdata(m_axi_rmem25___Stream2Mmap_25___mmap_RDATA),
    .s01_axi_rid(m_axi_rmem25___Stream2Mmap_25___mmap_RID),
    .s01_axi_rlast(m_axi_rmem25___Stream2Mmap_25___mmap_RLAST),
    .s01_axi_rready(m_axi_rmem25___Stream2Mmap_25___mmap_RREADY),
    .s01_axi_rresp(m_axi_rmem25___Stream2Mmap_25___mmap_RRESP),
    .s01_axi_rvalid(m_axi_rmem25___Stream2Mmap_25___mmap_RVALID),
    .s01_axi_wdata(m_axi_rmem25___Stream2Mmap_25___mmap_WDATA),
    .s01_axi_wlast(m_axi_rmem25___Stream2Mmap_25___mmap_WLAST),
    .s01_axi_wready(m_axi_rmem25___Stream2Mmap_25___mmap_WREADY),
    .s01_axi_wstrb(m_axi_rmem25___Stream2Mmap_25___mmap_WSTRB),
    .s01_axi_wvalid(m_axi_rmem25___Stream2Mmap_25___mmap_WVALID)
  );


  (* keep_hierarchy = "yes" *) axi_crossbar_2x1
  #(
    .DATA_WIDTH(512),
    .ADDR_WIDTH(64),
    .S_ID_WIDTH(1),
    .M_ID_WIDTH(2),
    .M00_ADDR_WIDTH(64),
    .M00_ISSUE(16),
    .S00_THREADS(1),
    .S01_THREADS(1)
  )
  axi_crossbar_2x1__rmem26
  (
    .clk(ap_clk),
    .rst(ap_rst_n_inv),
    .m00_axi_araddr(m_axi_rmem26_ARADDR),
    .m00_axi_arburst(m_axi_rmem26_ARBURST),
    .m00_axi_arcache(m_axi_rmem26_ARCACHE),
    .m00_axi_arid(m_axi_rmem26_ARID),
    .m00_axi_arlen(m_axi_rmem26_ARLEN),
    .m00_axi_arlock(m_axi_rmem26_ARLOCK),
    .m00_axi_arprot(m_axi_rmem26_ARPROT),
    .m00_axi_arqos(m_axi_rmem26_ARQOS),
    .m00_axi_arready(m_axi_rmem26_ARREADY),
    .m00_axi_arsize(m_axi_rmem26_ARSIZE),
    .m00_axi_arvalid(m_axi_rmem26_ARVALID),
    .m00_axi_awaddr(m_axi_rmem26_AWADDR),
    .m00_axi_awburst(m_axi_rmem26_AWBURST),
    .m00_axi_awcache(m_axi_rmem26_AWCACHE),
    .m00_axi_awid(m_axi_rmem26_AWID),
    .m00_axi_awlen(m_axi_rmem26_AWLEN),
    .m00_axi_awlock(m_axi_rmem26_AWLOCK),
    .m00_axi_awprot(m_axi_rmem26_AWPROT),
    .m00_axi_awqos(m_axi_rmem26_AWQOS),
    .m00_axi_awready(m_axi_rmem26_AWREADY),
    .m00_axi_awsize(m_axi_rmem26_AWSIZE),
    .m00_axi_awvalid(m_axi_rmem26_AWVALID),
    .m00_axi_bid(m_axi_rmem26_BID),
    .m00_axi_bready(m_axi_rmem26_BREADY),
    .m00_axi_bresp(m_axi_rmem26_BRESP),
    .m00_axi_bvalid(m_axi_rmem26_BVALID),
    .m00_axi_rdata(m_axi_rmem26_RDATA),
    .m00_axi_rid(m_axi_rmem26_RID),
    .m00_axi_rlast(m_axi_rmem26_RLAST),
    .m00_axi_rready(m_axi_rmem26_RREADY),
    .m00_axi_rresp(m_axi_rmem26_RRESP),
    .m00_axi_rvalid(m_axi_rmem26_RVALID),
    .m00_axi_wdata(m_axi_rmem26_WDATA),
    .m00_axi_wlast(m_axi_rmem26_WLAST),
    .m00_axi_wready(m_axi_rmem26_WREADY),
    .m00_axi_wstrb(m_axi_rmem26_WSTRB),
    .m00_axi_wvalid(m_axi_rmem26_WVALID),
    .s00_axi_araddr(m_axi_rmem26___Mmap2Stream_26___mmap_ARADDR),
    .s00_axi_arburst(m_axi_rmem26___Mmap2Stream_26___mmap_ARBURST),
    .s00_axi_arcache(m_axi_rmem26___Mmap2Stream_26___mmap_ARCACHE),
    .s00_axi_arid(m_axi_rmem26___Mmap2Stream_26___mmap_ARID),
    .s00_axi_arlen(m_axi_rmem26___Mmap2Stream_26___mmap_ARLEN),
    .s00_axi_arlock(m_axi_rmem26___Mmap2Stream_26___mmap_ARLOCK),
    .s00_axi_arprot(m_axi_rmem26___Mmap2Stream_26___mmap_ARPROT),
    .s00_axi_arqos(m_axi_rmem26___Mmap2Stream_26___mmap_ARQOS),
    .s00_axi_arready(m_axi_rmem26___Mmap2Stream_26___mmap_ARREADY),
    .s00_axi_arsize(m_axi_rmem26___Mmap2Stream_26___mmap_ARSIZE),
    .s00_axi_arvalid(m_axi_rmem26___Mmap2Stream_26___mmap_ARVALID),
    .s00_axi_awaddr(m_axi_rmem26___Mmap2Stream_26___mmap_AWADDR),
    .s00_axi_awburst(m_axi_rmem26___Mmap2Stream_26___mmap_AWBURST),
    .s00_axi_awcache(m_axi_rmem26___Mmap2Stream_26___mmap_AWCACHE),
    .s00_axi_awid(m_axi_rmem26___Mmap2Stream_26___mmap_AWID),
    .s00_axi_awlen(m_axi_rmem26___Mmap2Stream_26___mmap_AWLEN),
    .s00_axi_awlock(m_axi_rmem26___Mmap2Stream_26___mmap_AWLOCK),
    .s00_axi_awprot(m_axi_rmem26___Mmap2Stream_26___mmap_AWPROT),
    .s00_axi_awqos(m_axi_rmem26___Mmap2Stream_26___mmap_AWQOS),
    .s00_axi_awready(m_axi_rmem26___Mmap2Stream_26___mmap_AWREADY),
    .s00_axi_awsize(m_axi_rmem26___Mmap2Stream_26___mmap_AWSIZE),
    .s00_axi_awvalid(m_axi_rmem26___Mmap2Stream_26___mmap_AWVALID),
    .s00_axi_bid(m_axi_rmem26___Mmap2Stream_26___mmap_BID),
    .s00_axi_bready(m_axi_rmem26___Mmap2Stream_26___mmap_BREADY),
    .s00_axi_bresp(m_axi_rmem26___Mmap2Stream_26___mmap_BRESP),
    .s00_axi_bvalid(m_axi_rmem26___Mmap2Stream_26___mmap_BVALID),
    .s00_axi_rdata(m_axi_rmem26___Mmap2Stream_26___mmap_RDATA),
    .s00_axi_rid(m_axi_rmem26___Mmap2Stream_26___mmap_RID),
    .s00_axi_rlast(m_axi_rmem26___Mmap2Stream_26___mmap_RLAST),
    .s00_axi_rready(m_axi_rmem26___Mmap2Stream_26___mmap_RREADY),
    .s00_axi_rresp(m_axi_rmem26___Mmap2Stream_26___mmap_RRESP),
    .s00_axi_rvalid(m_axi_rmem26___Mmap2Stream_26___mmap_RVALID),
    .s00_axi_wdata(m_axi_rmem26___Mmap2Stream_26___mmap_WDATA),
    .s00_axi_wlast(m_axi_rmem26___Mmap2Stream_26___mmap_WLAST),
    .s00_axi_wready(m_axi_rmem26___Mmap2Stream_26___mmap_WREADY),
    .s00_axi_wstrb(m_axi_rmem26___Mmap2Stream_26___mmap_WSTRB),
    .s00_axi_wvalid(m_axi_rmem26___Mmap2Stream_26___mmap_WVALID),
    .s01_axi_araddr(m_axi_rmem26___Stream2Mmap_26___mmap_ARADDR),
    .s01_axi_arburst(m_axi_rmem26___Stream2Mmap_26___mmap_ARBURST),
    .s01_axi_arcache(m_axi_rmem26___Stream2Mmap_26___mmap_ARCACHE),
    .s01_axi_arid(m_axi_rmem26___Stream2Mmap_26___mmap_ARID),
    .s01_axi_arlen(m_axi_rmem26___Stream2Mmap_26___mmap_ARLEN),
    .s01_axi_arlock(m_axi_rmem26___Stream2Mmap_26___mmap_ARLOCK),
    .s01_axi_arprot(m_axi_rmem26___Stream2Mmap_26___mmap_ARPROT),
    .s01_axi_arqos(m_axi_rmem26___Stream2Mmap_26___mmap_ARQOS),
    .s01_axi_arready(m_axi_rmem26___Stream2Mmap_26___mmap_ARREADY),
    .s01_axi_arsize(m_axi_rmem26___Stream2Mmap_26___mmap_ARSIZE),
    .s01_axi_arvalid(m_axi_rmem26___Stream2Mmap_26___mmap_ARVALID),
    .s01_axi_awaddr(m_axi_rmem26___Stream2Mmap_26___mmap_AWADDR),
    .s01_axi_awburst(m_axi_rmem26___Stream2Mmap_26___mmap_AWBURST),
    .s01_axi_awcache(m_axi_rmem26___Stream2Mmap_26___mmap_AWCACHE),
    .s01_axi_awid(m_axi_rmem26___Stream2Mmap_26___mmap_AWID),
    .s01_axi_awlen(m_axi_rmem26___Stream2Mmap_26___mmap_AWLEN),
    .s01_axi_awlock(m_axi_rmem26___Stream2Mmap_26___mmap_AWLOCK),
    .s01_axi_awprot(m_axi_rmem26___Stream2Mmap_26___mmap_AWPROT),
    .s01_axi_awqos(m_axi_rmem26___Stream2Mmap_26___mmap_AWQOS),
    .s01_axi_awready(m_axi_rmem26___Stream2Mmap_26___mmap_AWREADY),
    .s01_axi_awsize(m_axi_rmem26___Stream2Mmap_26___mmap_AWSIZE),
    .s01_axi_awvalid(m_axi_rmem26___Stream2Mmap_26___mmap_AWVALID),
    .s01_axi_bid(m_axi_rmem26___Stream2Mmap_26___mmap_BID),
    .s01_axi_bready(m_axi_rmem26___Stream2Mmap_26___mmap_BREADY),
    .s01_axi_bresp(m_axi_rmem26___Stream2Mmap_26___mmap_BRESP),
    .s01_axi_bvalid(m_axi_rmem26___Stream2Mmap_26___mmap_BVALID),
    .s01_axi_rdata(m_axi_rmem26___Stream2Mmap_26___mmap_RDATA),
    .s01_axi_rid(m_axi_rmem26___Stream2Mmap_26___mmap_RID),
    .s01_axi_rlast(m_axi_rmem26___Stream2Mmap_26___mmap_RLAST),
    .s01_axi_rready(m_axi_rmem26___Stream2Mmap_26___mmap_RREADY),
    .s01_axi_rresp(m_axi_rmem26___Stream2Mmap_26___mmap_RRESP),
    .s01_axi_rvalid(m_axi_rmem26___Stream2Mmap_26___mmap_RVALID),
    .s01_axi_wdata(m_axi_rmem26___Stream2Mmap_26___mmap_WDATA),
    .s01_axi_wlast(m_axi_rmem26___Stream2Mmap_26___mmap_WLAST),
    .s01_axi_wready(m_axi_rmem26___Stream2Mmap_26___mmap_WREADY),
    .s01_axi_wstrb(m_axi_rmem26___Stream2Mmap_26___mmap_WSTRB),
    .s01_axi_wvalid(m_axi_rmem26___Stream2Mmap_26___mmap_WVALID)
  );


  (* keep_hierarchy = "yes" *) axi_crossbar_2x1
  #(
    .DATA_WIDTH(512),
    .ADDR_WIDTH(64),
    .S_ID_WIDTH(1),
    .M_ID_WIDTH(2),
    .M00_ADDR_WIDTH(64),
    .M00_ISSUE(16),
    .S00_THREADS(1),
    .S01_THREADS(1)
  )
  axi_crossbar_2x1__rmem27
  (
    .clk(ap_clk),
    .rst(ap_rst_n_inv),
    .m00_axi_araddr(m_axi_rmem27_ARADDR),
    .m00_axi_arburst(m_axi_rmem27_ARBURST),
    .m00_axi_arcache(m_axi_rmem27_ARCACHE),
    .m00_axi_arid(m_axi_rmem27_ARID),
    .m00_axi_arlen(m_axi_rmem27_ARLEN),
    .m00_axi_arlock(m_axi_rmem27_ARLOCK),
    .m00_axi_arprot(m_axi_rmem27_ARPROT),
    .m00_axi_arqos(m_axi_rmem27_ARQOS),
    .m00_axi_arready(m_axi_rmem27_ARREADY),
    .m00_axi_arsize(m_axi_rmem27_ARSIZE),
    .m00_axi_arvalid(m_axi_rmem27_ARVALID),
    .m00_axi_awaddr(m_axi_rmem27_AWADDR),
    .m00_axi_awburst(m_axi_rmem27_AWBURST),
    .m00_axi_awcache(m_axi_rmem27_AWCACHE),
    .m00_axi_awid(m_axi_rmem27_AWID),
    .m00_axi_awlen(m_axi_rmem27_AWLEN),
    .m00_axi_awlock(m_axi_rmem27_AWLOCK),
    .m00_axi_awprot(m_axi_rmem27_AWPROT),
    .m00_axi_awqos(m_axi_rmem27_AWQOS),
    .m00_axi_awready(m_axi_rmem27_AWREADY),
    .m00_axi_awsize(m_axi_rmem27_AWSIZE),
    .m00_axi_awvalid(m_axi_rmem27_AWVALID),
    .m00_axi_bid(m_axi_rmem27_BID),
    .m00_axi_bready(m_axi_rmem27_BREADY),
    .m00_axi_bresp(m_axi_rmem27_BRESP),
    .m00_axi_bvalid(m_axi_rmem27_BVALID),
    .m00_axi_rdata(m_axi_rmem27_RDATA),
    .m00_axi_rid(m_axi_rmem27_RID),
    .m00_axi_rlast(m_axi_rmem27_RLAST),
    .m00_axi_rready(m_axi_rmem27_RREADY),
    .m00_axi_rresp(m_axi_rmem27_RRESP),
    .m00_axi_rvalid(m_axi_rmem27_RVALID),
    .m00_axi_wdata(m_axi_rmem27_WDATA),
    .m00_axi_wlast(m_axi_rmem27_WLAST),
    .m00_axi_wready(m_axi_rmem27_WREADY),
    .m00_axi_wstrb(m_axi_rmem27_WSTRB),
    .m00_axi_wvalid(m_axi_rmem27_WVALID),
    .s00_axi_araddr(m_axi_rmem27___Mmap2Stream_27___mmap_ARADDR),
    .s00_axi_arburst(m_axi_rmem27___Mmap2Stream_27___mmap_ARBURST),
    .s00_axi_arcache(m_axi_rmem27___Mmap2Stream_27___mmap_ARCACHE),
    .s00_axi_arid(m_axi_rmem27___Mmap2Stream_27___mmap_ARID),
    .s00_axi_arlen(m_axi_rmem27___Mmap2Stream_27___mmap_ARLEN),
    .s00_axi_arlock(m_axi_rmem27___Mmap2Stream_27___mmap_ARLOCK),
    .s00_axi_arprot(m_axi_rmem27___Mmap2Stream_27___mmap_ARPROT),
    .s00_axi_arqos(m_axi_rmem27___Mmap2Stream_27___mmap_ARQOS),
    .s00_axi_arready(m_axi_rmem27___Mmap2Stream_27___mmap_ARREADY),
    .s00_axi_arsize(m_axi_rmem27___Mmap2Stream_27___mmap_ARSIZE),
    .s00_axi_arvalid(m_axi_rmem27___Mmap2Stream_27___mmap_ARVALID),
    .s00_axi_awaddr(m_axi_rmem27___Mmap2Stream_27___mmap_AWADDR),
    .s00_axi_awburst(m_axi_rmem27___Mmap2Stream_27___mmap_AWBURST),
    .s00_axi_awcache(m_axi_rmem27___Mmap2Stream_27___mmap_AWCACHE),
    .s00_axi_awid(m_axi_rmem27___Mmap2Stream_27___mmap_AWID),
    .s00_axi_awlen(m_axi_rmem27___Mmap2Stream_27___mmap_AWLEN),
    .s00_axi_awlock(m_axi_rmem27___Mmap2Stream_27___mmap_AWLOCK),
    .s00_axi_awprot(m_axi_rmem27___Mmap2Stream_27___mmap_AWPROT),
    .s00_axi_awqos(m_axi_rmem27___Mmap2Stream_27___mmap_AWQOS),
    .s00_axi_awready(m_axi_rmem27___Mmap2Stream_27___mmap_AWREADY),
    .s00_axi_awsize(m_axi_rmem27___Mmap2Stream_27___mmap_AWSIZE),
    .s00_axi_awvalid(m_axi_rmem27___Mmap2Stream_27___mmap_AWVALID),
    .s00_axi_bid(m_axi_rmem27___Mmap2Stream_27___mmap_BID),
    .s00_axi_bready(m_axi_rmem27___Mmap2Stream_27___mmap_BREADY),
    .s00_axi_bresp(m_axi_rmem27___Mmap2Stream_27___mmap_BRESP),
    .s00_axi_bvalid(m_axi_rmem27___Mmap2Stream_27___mmap_BVALID),
    .s00_axi_rdata(m_axi_rmem27___Mmap2Stream_27___mmap_RDATA),
    .s00_axi_rid(m_axi_rmem27___Mmap2Stream_27___mmap_RID),
    .s00_axi_rlast(m_axi_rmem27___Mmap2Stream_27___mmap_RLAST),
    .s00_axi_rready(m_axi_rmem27___Mmap2Stream_27___mmap_RREADY),
    .s00_axi_rresp(m_axi_rmem27___Mmap2Stream_27___mmap_RRESP),
    .s00_axi_rvalid(m_axi_rmem27___Mmap2Stream_27___mmap_RVALID),
    .s00_axi_wdata(m_axi_rmem27___Mmap2Stream_27___mmap_WDATA),
    .s00_axi_wlast(m_axi_rmem27___Mmap2Stream_27___mmap_WLAST),
    .s00_axi_wready(m_axi_rmem27___Mmap2Stream_27___mmap_WREADY),
    .s00_axi_wstrb(m_axi_rmem27___Mmap2Stream_27___mmap_WSTRB),
    .s00_axi_wvalid(m_axi_rmem27___Mmap2Stream_27___mmap_WVALID),
    .s01_axi_araddr(m_axi_rmem27___Stream2Mmap_27___mmap_ARADDR),
    .s01_axi_arburst(m_axi_rmem27___Stream2Mmap_27___mmap_ARBURST),
    .s01_axi_arcache(m_axi_rmem27___Stream2Mmap_27___mmap_ARCACHE),
    .s01_axi_arid(m_axi_rmem27___Stream2Mmap_27___mmap_ARID),
    .s01_axi_arlen(m_axi_rmem27___Stream2Mmap_27___mmap_ARLEN),
    .s01_axi_arlock(m_axi_rmem27___Stream2Mmap_27___mmap_ARLOCK),
    .s01_axi_arprot(m_axi_rmem27___Stream2Mmap_27___mmap_ARPROT),
    .s01_axi_arqos(m_axi_rmem27___Stream2Mmap_27___mmap_ARQOS),
    .s01_axi_arready(m_axi_rmem27___Stream2Mmap_27___mmap_ARREADY),
    .s01_axi_arsize(m_axi_rmem27___Stream2Mmap_27___mmap_ARSIZE),
    .s01_axi_arvalid(m_axi_rmem27___Stream2Mmap_27___mmap_ARVALID),
    .s01_axi_awaddr(m_axi_rmem27___Stream2Mmap_27___mmap_AWADDR),
    .s01_axi_awburst(m_axi_rmem27___Stream2Mmap_27___mmap_AWBURST),
    .s01_axi_awcache(m_axi_rmem27___Stream2Mmap_27___mmap_AWCACHE),
    .s01_axi_awid(m_axi_rmem27___Stream2Mmap_27___mmap_AWID),
    .s01_axi_awlen(m_axi_rmem27___Stream2Mmap_27___mmap_AWLEN),
    .s01_axi_awlock(m_axi_rmem27___Stream2Mmap_27___mmap_AWLOCK),
    .s01_axi_awprot(m_axi_rmem27___Stream2Mmap_27___mmap_AWPROT),
    .s01_axi_awqos(m_axi_rmem27___Stream2Mmap_27___mmap_AWQOS),
    .s01_axi_awready(m_axi_rmem27___Stream2Mmap_27___mmap_AWREADY),
    .s01_axi_awsize(m_axi_rmem27___Stream2Mmap_27___mmap_AWSIZE),
    .s01_axi_awvalid(m_axi_rmem27___Stream2Mmap_27___mmap_AWVALID),
    .s01_axi_bid(m_axi_rmem27___Stream2Mmap_27___mmap_BID),
    .s01_axi_bready(m_axi_rmem27___Stream2Mmap_27___mmap_BREADY),
    .s01_axi_bresp(m_axi_rmem27___Stream2Mmap_27___mmap_BRESP),
    .s01_axi_bvalid(m_axi_rmem27___Stream2Mmap_27___mmap_BVALID),
    .s01_axi_rdata(m_axi_rmem27___Stream2Mmap_27___mmap_RDATA),
    .s01_axi_rid(m_axi_rmem27___Stream2Mmap_27___mmap_RID),
    .s01_axi_rlast(m_axi_rmem27___Stream2Mmap_27___mmap_RLAST),
    .s01_axi_rready(m_axi_rmem27___Stream2Mmap_27___mmap_RREADY),
    .s01_axi_rresp(m_axi_rmem27___Stream2Mmap_27___mmap_RRESP),
    .s01_axi_rvalid(m_axi_rmem27___Stream2Mmap_27___mmap_RVALID),
    .s01_axi_wdata(m_axi_rmem27___Stream2Mmap_27___mmap_WDATA),
    .s01_axi_wlast(m_axi_rmem27___Stream2Mmap_27___mmap_WLAST),
    .s01_axi_wready(m_axi_rmem27___Stream2Mmap_27___mmap_WREADY),
    .s01_axi_wstrb(m_axi_rmem27___Stream2Mmap_27___mmap_WSTRB),
    .s01_axi_wvalid(m_axi_rmem27___Stream2Mmap_27___mmap_WVALID)
  );


  (* keep_hierarchy = "yes" *) Mmap2Stream
  Mmap2Stream_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Mmap2Stream_0__ap_start),
    .ap_done(Mmap2Stream_0__ap_done),
    .ap_idle(Mmap2Stream_0__ap_idle),
    .ap_ready(Mmap2Stream_0__ap_ready),
    .n(Mmap2Stream_0___n__q0),
    .stream_din(qr0_vadd_bw__din),
    .stream_full_n(qr0_vadd_bw__full_n),
    .stream_write(qr0_vadd_bw__write),
    .m_axi_mmap_ARADDR(m_axi_rmem0___Mmap2Stream_0___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem0___Mmap2Stream_0___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem0___Mmap2Stream_0___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem0___Mmap2Stream_0___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem0___Mmap2Stream_0___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem0___Mmap2Stream_0___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem0___Mmap2Stream_0___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem0___Mmap2Stream_0___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem0___Mmap2Stream_0___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem0___Mmap2Stream_0___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem0___Mmap2Stream_0___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem0___Mmap2Stream_0___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem0___Mmap2Stream_0___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem0___Mmap2Stream_0___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem0___Mmap2Stream_0___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem0___Mmap2Stream_0___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem0___Mmap2Stream_0___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem0___Mmap2Stream_0___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem0___Mmap2Stream_0___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem0___Mmap2Stream_0___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem0___Mmap2Stream_0___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem0___Mmap2Stream_0___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem0___Mmap2Stream_0___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem0___Mmap2Stream_0___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem0___Mmap2Stream_0___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem0___Mmap2Stream_0___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem0___Mmap2Stream_0___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem0___Mmap2Stream_0___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem0___Mmap2Stream_0___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem0___Mmap2Stream_0___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem0___Mmap2Stream_0___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem0___Mmap2Stream_0___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem0___Mmap2Stream_0___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem0___Mmap2Stream_0___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem0___Mmap2Stream_0___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem0___Mmap2Stream_0___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem0___Mmap2Stream_0___mmap_AWQOS),
    .mmap_offset(Mmap2Stream_0___rmem0__q0)
  );


  (* keep_hierarchy = "yes" *) Mmap2Stream
  Mmap2Stream_1
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Mmap2Stream_1__ap_start),
    .ap_done(Mmap2Stream_1__ap_done),
    .ap_idle(Mmap2Stream_1__ap_idle),
    .ap_ready(Mmap2Stream_1__ap_ready),
    .n(Mmap2Stream_1___n__q0),
    .stream_din(qr1_vadd_bw__din),
    .stream_full_n(qr1_vadd_bw__full_n),
    .stream_write(qr1_vadd_bw__write),
    .m_axi_mmap_ARADDR(m_axi_rmem1___Mmap2Stream_1___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem1___Mmap2Stream_1___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem1___Mmap2Stream_1___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem1___Mmap2Stream_1___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem1___Mmap2Stream_1___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem1___Mmap2Stream_1___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem1___Mmap2Stream_1___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem1___Mmap2Stream_1___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem1___Mmap2Stream_1___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem1___Mmap2Stream_1___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem1___Mmap2Stream_1___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem1___Mmap2Stream_1___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem1___Mmap2Stream_1___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem1___Mmap2Stream_1___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem1___Mmap2Stream_1___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem1___Mmap2Stream_1___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem1___Mmap2Stream_1___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem1___Mmap2Stream_1___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem1___Mmap2Stream_1___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem1___Mmap2Stream_1___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem1___Mmap2Stream_1___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem1___Mmap2Stream_1___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem1___Mmap2Stream_1___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem1___Mmap2Stream_1___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem1___Mmap2Stream_1___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem1___Mmap2Stream_1___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem1___Mmap2Stream_1___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem1___Mmap2Stream_1___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem1___Mmap2Stream_1___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem1___Mmap2Stream_1___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem1___Mmap2Stream_1___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem1___Mmap2Stream_1___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem1___Mmap2Stream_1___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem1___Mmap2Stream_1___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem1___Mmap2Stream_1___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem1___Mmap2Stream_1___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem1___Mmap2Stream_1___mmap_AWQOS),
    .mmap_offset(Mmap2Stream_1___rmem1__q0)
  );


  (* keep_hierarchy = "yes" *) Mmap2Stream
  Mmap2Stream_2
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Mmap2Stream_2__ap_start),
    .ap_done(Mmap2Stream_2__ap_done),
    .ap_idle(Mmap2Stream_2__ap_idle),
    .ap_ready(Mmap2Stream_2__ap_ready),
    .n(Mmap2Stream_2___n__q0),
    .stream_din(qr2_vadd_bw__din),
    .stream_full_n(qr2_vadd_bw__full_n),
    .stream_write(qr2_vadd_bw__write),
    .m_axi_mmap_ARADDR(m_axi_rmem2___Mmap2Stream_2___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem2___Mmap2Stream_2___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem2___Mmap2Stream_2___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem2___Mmap2Stream_2___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem2___Mmap2Stream_2___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem2___Mmap2Stream_2___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem2___Mmap2Stream_2___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem2___Mmap2Stream_2___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem2___Mmap2Stream_2___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem2___Mmap2Stream_2___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem2___Mmap2Stream_2___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem2___Mmap2Stream_2___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem2___Mmap2Stream_2___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem2___Mmap2Stream_2___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem2___Mmap2Stream_2___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem2___Mmap2Stream_2___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem2___Mmap2Stream_2___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem2___Mmap2Stream_2___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem2___Mmap2Stream_2___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem2___Mmap2Stream_2___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem2___Mmap2Stream_2___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem2___Mmap2Stream_2___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem2___Mmap2Stream_2___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem2___Mmap2Stream_2___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem2___Mmap2Stream_2___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem2___Mmap2Stream_2___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem2___Mmap2Stream_2___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem2___Mmap2Stream_2___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem2___Mmap2Stream_2___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem2___Mmap2Stream_2___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem2___Mmap2Stream_2___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem2___Mmap2Stream_2___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem2___Mmap2Stream_2___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem2___Mmap2Stream_2___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem2___Mmap2Stream_2___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem2___Mmap2Stream_2___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem2___Mmap2Stream_2___mmap_AWQOS),
    .mmap_offset(Mmap2Stream_2___rmem2__q0)
  );


  (* keep_hierarchy = "yes" *) Mmap2Stream
  Mmap2Stream_3
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Mmap2Stream_3__ap_start),
    .ap_done(Mmap2Stream_3__ap_done),
    .ap_idle(Mmap2Stream_3__ap_idle),
    .ap_ready(Mmap2Stream_3__ap_ready),
    .n(Mmap2Stream_3___n__q0),
    .stream_din(qr3_vadd_bw__din),
    .stream_full_n(qr3_vadd_bw__full_n),
    .stream_write(qr3_vadd_bw__write),
    .m_axi_mmap_ARADDR(m_axi_rmem3___Mmap2Stream_3___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem3___Mmap2Stream_3___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem3___Mmap2Stream_3___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem3___Mmap2Stream_3___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem3___Mmap2Stream_3___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem3___Mmap2Stream_3___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem3___Mmap2Stream_3___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem3___Mmap2Stream_3___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem3___Mmap2Stream_3___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem3___Mmap2Stream_3___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem3___Mmap2Stream_3___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem3___Mmap2Stream_3___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem3___Mmap2Stream_3___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem3___Mmap2Stream_3___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem3___Mmap2Stream_3___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem3___Mmap2Stream_3___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem3___Mmap2Stream_3___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem3___Mmap2Stream_3___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem3___Mmap2Stream_3___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem3___Mmap2Stream_3___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem3___Mmap2Stream_3___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem3___Mmap2Stream_3___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem3___Mmap2Stream_3___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem3___Mmap2Stream_3___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem3___Mmap2Stream_3___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem3___Mmap2Stream_3___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem3___Mmap2Stream_3___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem3___Mmap2Stream_3___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem3___Mmap2Stream_3___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem3___Mmap2Stream_3___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem3___Mmap2Stream_3___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem3___Mmap2Stream_3___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem3___Mmap2Stream_3___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem3___Mmap2Stream_3___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem3___Mmap2Stream_3___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem3___Mmap2Stream_3___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem3___Mmap2Stream_3___mmap_AWQOS),
    .mmap_offset(Mmap2Stream_3___rmem3__q0)
  );


  (* keep_hierarchy = "yes" *) Mmap2Stream
  Mmap2Stream_4
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Mmap2Stream_4__ap_start),
    .ap_done(Mmap2Stream_4__ap_done),
    .ap_idle(Mmap2Stream_4__ap_idle),
    .ap_ready(Mmap2Stream_4__ap_ready),
    .n(Mmap2Stream_4___n__q0),
    .stream_din(qr4_vadd_bw__din),
    .stream_full_n(qr4_vadd_bw__full_n),
    .stream_write(qr4_vadd_bw__write),
    .m_axi_mmap_ARADDR(m_axi_rmem4___Mmap2Stream_4___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem4___Mmap2Stream_4___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem4___Mmap2Stream_4___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem4___Mmap2Stream_4___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem4___Mmap2Stream_4___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem4___Mmap2Stream_4___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem4___Mmap2Stream_4___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem4___Mmap2Stream_4___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem4___Mmap2Stream_4___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem4___Mmap2Stream_4___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem4___Mmap2Stream_4___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem4___Mmap2Stream_4___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem4___Mmap2Stream_4___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem4___Mmap2Stream_4___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem4___Mmap2Stream_4___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem4___Mmap2Stream_4___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem4___Mmap2Stream_4___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem4___Mmap2Stream_4___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem4___Mmap2Stream_4___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem4___Mmap2Stream_4___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem4___Mmap2Stream_4___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem4___Mmap2Stream_4___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem4___Mmap2Stream_4___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem4___Mmap2Stream_4___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem4___Mmap2Stream_4___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem4___Mmap2Stream_4___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem4___Mmap2Stream_4___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem4___Mmap2Stream_4___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem4___Mmap2Stream_4___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem4___Mmap2Stream_4___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem4___Mmap2Stream_4___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem4___Mmap2Stream_4___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem4___Mmap2Stream_4___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem4___Mmap2Stream_4___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem4___Mmap2Stream_4___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem4___Mmap2Stream_4___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem4___Mmap2Stream_4___mmap_AWQOS),
    .mmap_offset(Mmap2Stream_4___rmem4__q0)
  );


  (* keep_hierarchy = "yes" *) Mmap2Stream
  Mmap2Stream_5
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Mmap2Stream_5__ap_start),
    .ap_done(Mmap2Stream_5__ap_done),
    .ap_idle(Mmap2Stream_5__ap_idle),
    .ap_ready(Mmap2Stream_5__ap_ready),
    .n(Mmap2Stream_5___n__q0),
    .stream_din(qr5_vadd_bw__din),
    .stream_full_n(qr5_vadd_bw__full_n),
    .stream_write(qr5_vadd_bw__write),
    .m_axi_mmap_ARADDR(m_axi_rmem5___Mmap2Stream_5___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem5___Mmap2Stream_5___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem5___Mmap2Stream_5___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem5___Mmap2Stream_5___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem5___Mmap2Stream_5___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem5___Mmap2Stream_5___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem5___Mmap2Stream_5___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem5___Mmap2Stream_5___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem5___Mmap2Stream_5___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem5___Mmap2Stream_5___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem5___Mmap2Stream_5___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem5___Mmap2Stream_5___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem5___Mmap2Stream_5___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem5___Mmap2Stream_5___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem5___Mmap2Stream_5___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem5___Mmap2Stream_5___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem5___Mmap2Stream_5___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem5___Mmap2Stream_5___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem5___Mmap2Stream_5___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem5___Mmap2Stream_5___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem5___Mmap2Stream_5___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem5___Mmap2Stream_5___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem5___Mmap2Stream_5___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem5___Mmap2Stream_5___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem5___Mmap2Stream_5___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem5___Mmap2Stream_5___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem5___Mmap2Stream_5___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem5___Mmap2Stream_5___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem5___Mmap2Stream_5___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem5___Mmap2Stream_5___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem5___Mmap2Stream_5___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem5___Mmap2Stream_5___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem5___Mmap2Stream_5___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem5___Mmap2Stream_5___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem5___Mmap2Stream_5___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem5___Mmap2Stream_5___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem5___Mmap2Stream_5___mmap_AWQOS),
    .mmap_offset(Mmap2Stream_5___rmem5__q0)
  );


  (* keep_hierarchy = "yes" *) Mmap2Stream
  Mmap2Stream_6
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Mmap2Stream_6__ap_start),
    .ap_done(Mmap2Stream_6__ap_done),
    .ap_idle(Mmap2Stream_6__ap_idle),
    .ap_ready(Mmap2Stream_6__ap_ready),
    .n(Mmap2Stream_6___n__q0),
    .stream_din(qr6_vadd_bw__din),
    .stream_full_n(qr6_vadd_bw__full_n),
    .stream_write(qr6_vadd_bw__write),
    .m_axi_mmap_ARADDR(m_axi_rmem6___Mmap2Stream_6___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem6___Mmap2Stream_6___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem6___Mmap2Stream_6___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem6___Mmap2Stream_6___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem6___Mmap2Stream_6___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem6___Mmap2Stream_6___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem6___Mmap2Stream_6___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem6___Mmap2Stream_6___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem6___Mmap2Stream_6___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem6___Mmap2Stream_6___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem6___Mmap2Stream_6___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem6___Mmap2Stream_6___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem6___Mmap2Stream_6___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem6___Mmap2Stream_6___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem6___Mmap2Stream_6___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem6___Mmap2Stream_6___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem6___Mmap2Stream_6___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem6___Mmap2Stream_6___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem6___Mmap2Stream_6___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem6___Mmap2Stream_6___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem6___Mmap2Stream_6___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem6___Mmap2Stream_6___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem6___Mmap2Stream_6___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem6___Mmap2Stream_6___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem6___Mmap2Stream_6___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem6___Mmap2Stream_6___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem6___Mmap2Stream_6___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem6___Mmap2Stream_6___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem6___Mmap2Stream_6___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem6___Mmap2Stream_6___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem6___Mmap2Stream_6___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem6___Mmap2Stream_6___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem6___Mmap2Stream_6___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem6___Mmap2Stream_6___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem6___Mmap2Stream_6___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem6___Mmap2Stream_6___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem6___Mmap2Stream_6___mmap_AWQOS),
    .mmap_offset(Mmap2Stream_6___rmem6__q0)
  );


  (* keep_hierarchy = "yes" *) Mmap2Stream
  Mmap2Stream_7
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Mmap2Stream_7__ap_start),
    .ap_done(Mmap2Stream_7__ap_done),
    .ap_idle(Mmap2Stream_7__ap_idle),
    .ap_ready(Mmap2Stream_7__ap_ready),
    .n(Mmap2Stream_7___n__q0),
    .stream_din(qr7_vadd_bw__din),
    .stream_full_n(qr7_vadd_bw__full_n),
    .stream_write(qr7_vadd_bw__write),
    .m_axi_mmap_ARADDR(m_axi_rmem7___Mmap2Stream_7___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem7___Mmap2Stream_7___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem7___Mmap2Stream_7___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem7___Mmap2Stream_7___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem7___Mmap2Stream_7___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem7___Mmap2Stream_7___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem7___Mmap2Stream_7___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem7___Mmap2Stream_7___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem7___Mmap2Stream_7___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem7___Mmap2Stream_7___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem7___Mmap2Stream_7___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem7___Mmap2Stream_7___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem7___Mmap2Stream_7___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem7___Mmap2Stream_7___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem7___Mmap2Stream_7___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem7___Mmap2Stream_7___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem7___Mmap2Stream_7___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem7___Mmap2Stream_7___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem7___Mmap2Stream_7___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem7___Mmap2Stream_7___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem7___Mmap2Stream_7___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem7___Mmap2Stream_7___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem7___Mmap2Stream_7___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem7___Mmap2Stream_7___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem7___Mmap2Stream_7___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem7___Mmap2Stream_7___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem7___Mmap2Stream_7___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem7___Mmap2Stream_7___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem7___Mmap2Stream_7___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem7___Mmap2Stream_7___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem7___Mmap2Stream_7___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem7___Mmap2Stream_7___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem7___Mmap2Stream_7___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem7___Mmap2Stream_7___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem7___Mmap2Stream_7___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem7___Mmap2Stream_7___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem7___Mmap2Stream_7___mmap_AWQOS),
    .mmap_offset(Mmap2Stream_7___rmem7__q0)
  );


  (* keep_hierarchy = "yes" *) Mmap2Stream
  Mmap2Stream_8
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Mmap2Stream_8__ap_start),
    .ap_done(Mmap2Stream_8__ap_done),
    .ap_idle(Mmap2Stream_8__ap_idle),
    .ap_ready(Mmap2Stream_8__ap_ready),
    .n(Mmap2Stream_8___n__q0),
    .stream_din(qr8_vadd_bw__din),
    .stream_full_n(qr8_vadd_bw__full_n),
    .stream_write(qr8_vadd_bw__write),
    .m_axi_mmap_ARADDR(m_axi_rmem8___Mmap2Stream_8___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem8___Mmap2Stream_8___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem8___Mmap2Stream_8___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem8___Mmap2Stream_8___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem8___Mmap2Stream_8___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem8___Mmap2Stream_8___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem8___Mmap2Stream_8___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem8___Mmap2Stream_8___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem8___Mmap2Stream_8___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem8___Mmap2Stream_8___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem8___Mmap2Stream_8___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem8___Mmap2Stream_8___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem8___Mmap2Stream_8___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem8___Mmap2Stream_8___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem8___Mmap2Stream_8___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem8___Mmap2Stream_8___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem8___Mmap2Stream_8___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem8___Mmap2Stream_8___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem8___Mmap2Stream_8___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem8___Mmap2Stream_8___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem8___Mmap2Stream_8___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem8___Mmap2Stream_8___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem8___Mmap2Stream_8___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem8___Mmap2Stream_8___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem8___Mmap2Stream_8___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem8___Mmap2Stream_8___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem8___Mmap2Stream_8___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem8___Mmap2Stream_8___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem8___Mmap2Stream_8___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem8___Mmap2Stream_8___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem8___Mmap2Stream_8___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem8___Mmap2Stream_8___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem8___Mmap2Stream_8___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem8___Mmap2Stream_8___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem8___Mmap2Stream_8___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem8___Mmap2Stream_8___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem8___Mmap2Stream_8___mmap_AWQOS),
    .mmap_offset(Mmap2Stream_8___rmem8__q0)
  );


  (* keep_hierarchy = "yes" *) Mmap2Stream
  Mmap2Stream_9
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Mmap2Stream_9__ap_start),
    .ap_done(Mmap2Stream_9__ap_done),
    .ap_idle(Mmap2Stream_9__ap_idle),
    .ap_ready(Mmap2Stream_9__ap_ready),
    .n(Mmap2Stream_9___n__q0),
    .stream_din(qr9_vadd_bw__din),
    .stream_full_n(qr9_vadd_bw__full_n),
    .stream_write(qr9_vadd_bw__write),
    .m_axi_mmap_ARADDR(m_axi_rmem9___Mmap2Stream_9___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem9___Mmap2Stream_9___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem9___Mmap2Stream_9___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem9___Mmap2Stream_9___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem9___Mmap2Stream_9___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem9___Mmap2Stream_9___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem9___Mmap2Stream_9___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem9___Mmap2Stream_9___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem9___Mmap2Stream_9___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem9___Mmap2Stream_9___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem9___Mmap2Stream_9___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem9___Mmap2Stream_9___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem9___Mmap2Stream_9___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem9___Mmap2Stream_9___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem9___Mmap2Stream_9___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem9___Mmap2Stream_9___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem9___Mmap2Stream_9___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem9___Mmap2Stream_9___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem9___Mmap2Stream_9___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem9___Mmap2Stream_9___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem9___Mmap2Stream_9___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem9___Mmap2Stream_9___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem9___Mmap2Stream_9___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem9___Mmap2Stream_9___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem9___Mmap2Stream_9___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem9___Mmap2Stream_9___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem9___Mmap2Stream_9___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem9___Mmap2Stream_9___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem9___Mmap2Stream_9___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem9___Mmap2Stream_9___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem9___Mmap2Stream_9___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem9___Mmap2Stream_9___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem9___Mmap2Stream_9___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem9___Mmap2Stream_9___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem9___Mmap2Stream_9___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem9___Mmap2Stream_9___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem9___Mmap2Stream_9___mmap_AWQOS),
    .mmap_offset(Mmap2Stream_9___rmem9__q0)
  );


  (* keep_hierarchy = "yes" *) Mmap2Stream
  Mmap2Stream_10
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Mmap2Stream_10__ap_start),
    .ap_done(Mmap2Stream_10__ap_done),
    .ap_idle(Mmap2Stream_10__ap_idle),
    .ap_ready(Mmap2Stream_10__ap_ready),
    .n(Mmap2Stream_10___n__q0),
    .stream_din(qr10_vadd_bw__din),
    .stream_full_n(qr10_vadd_bw__full_n),
    .stream_write(qr10_vadd_bw__write),
    .m_axi_mmap_ARADDR(m_axi_rmem10___Mmap2Stream_10___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem10___Mmap2Stream_10___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem10___Mmap2Stream_10___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem10___Mmap2Stream_10___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem10___Mmap2Stream_10___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem10___Mmap2Stream_10___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem10___Mmap2Stream_10___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem10___Mmap2Stream_10___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem10___Mmap2Stream_10___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem10___Mmap2Stream_10___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem10___Mmap2Stream_10___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem10___Mmap2Stream_10___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem10___Mmap2Stream_10___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem10___Mmap2Stream_10___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem10___Mmap2Stream_10___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem10___Mmap2Stream_10___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem10___Mmap2Stream_10___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem10___Mmap2Stream_10___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem10___Mmap2Stream_10___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem10___Mmap2Stream_10___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem10___Mmap2Stream_10___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem10___Mmap2Stream_10___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem10___Mmap2Stream_10___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem10___Mmap2Stream_10___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem10___Mmap2Stream_10___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem10___Mmap2Stream_10___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem10___Mmap2Stream_10___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem10___Mmap2Stream_10___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem10___Mmap2Stream_10___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem10___Mmap2Stream_10___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem10___Mmap2Stream_10___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem10___Mmap2Stream_10___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem10___Mmap2Stream_10___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem10___Mmap2Stream_10___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem10___Mmap2Stream_10___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem10___Mmap2Stream_10___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem10___Mmap2Stream_10___mmap_AWQOS),
    .mmap_offset(Mmap2Stream_10___rmem10__q0)
  );


  (* keep_hierarchy = "yes" *) Mmap2Stream
  Mmap2Stream_11
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Mmap2Stream_11__ap_start),
    .ap_done(Mmap2Stream_11__ap_done),
    .ap_idle(Mmap2Stream_11__ap_idle),
    .ap_ready(Mmap2Stream_11__ap_ready),
    .n(Mmap2Stream_11___n__q0),
    .stream_din(qr11_vadd_bw__din),
    .stream_full_n(qr11_vadd_bw__full_n),
    .stream_write(qr11_vadd_bw__write),
    .m_axi_mmap_ARADDR(m_axi_rmem11___Mmap2Stream_11___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem11___Mmap2Stream_11___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem11___Mmap2Stream_11___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem11___Mmap2Stream_11___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem11___Mmap2Stream_11___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem11___Mmap2Stream_11___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem11___Mmap2Stream_11___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem11___Mmap2Stream_11___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem11___Mmap2Stream_11___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem11___Mmap2Stream_11___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem11___Mmap2Stream_11___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem11___Mmap2Stream_11___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem11___Mmap2Stream_11___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem11___Mmap2Stream_11___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem11___Mmap2Stream_11___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem11___Mmap2Stream_11___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem11___Mmap2Stream_11___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem11___Mmap2Stream_11___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem11___Mmap2Stream_11___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem11___Mmap2Stream_11___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem11___Mmap2Stream_11___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem11___Mmap2Stream_11___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem11___Mmap2Stream_11___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem11___Mmap2Stream_11___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem11___Mmap2Stream_11___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem11___Mmap2Stream_11___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem11___Mmap2Stream_11___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem11___Mmap2Stream_11___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem11___Mmap2Stream_11___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem11___Mmap2Stream_11___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem11___Mmap2Stream_11___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem11___Mmap2Stream_11___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem11___Mmap2Stream_11___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem11___Mmap2Stream_11___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem11___Mmap2Stream_11___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem11___Mmap2Stream_11___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem11___Mmap2Stream_11___mmap_AWQOS),
    .mmap_offset(Mmap2Stream_11___rmem11__q0)
  );


  (* keep_hierarchy = "yes" *) Mmap2Stream
  Mmap2Stream_12
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Mmap2Stream_12__ap_start),
    .ap_done(Mmap2Stream_12__ap_done),
    .ap_idle(Mmap2Stream_12__ap_idle),
    .ap_ready(Mmap2Stream_12__ap_ready),
    .n(Mmap2Stream_12___n__q0),
    .stream_din(qr12_vadd_bw__din),
    .stream_full_n(qr12_vadd_bw__full_n),
    .stream_write(qr12_vadd_bw__write),
    .m_axi_mmap_ARADDR(m_axi_rmem12___Mmap2Stream_12___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem12___Mmap2Stream_12___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem12___Mmap2Stream_12___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem12___Mmap2Stream_12___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem12___Mmap2Stream_12___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem12___Mmap2Stream_12___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem12___Mmap2Stream_12___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem12___Mmap2Stream_12___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem12___Mmap2Stream_12___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem12___Mmap2Stream_12___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem12___Mmap2Stream_12___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem12___Mmap2Stream_12___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem12___Mmap2Stream_12___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem12___Mmap2Stream_12___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem12___Mmap2Stream_12___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem12___Mmap2Stream_12___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem12___Mmap2Stream_12___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem12___Mmap2Stream_12___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem12___Mmap2Stream_12___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem12___Mmap2Stream_12___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem12___Mmap2Stream_12___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem12___Mmap2Stream_12___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem12___Mmap2Stream_12___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem12___Mmap2Stream_12___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem12___Mmap2Stream_12___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem12___Mmap2Stream_12___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem12___Mmap2Stream_12___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem12___Mmap2Stream_12___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem12___Mmap2Stream_12___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem12___Mmap2Stream_12___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem12___Mmap2Stream_12___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem12___Mmap2Stream_12___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem12___Mmap2Stream_12___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem12___Mmap2Stream_12___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem12___Mmap2Stream_12___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem12___Mmap2Stream_12___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem12___Mmap2Stream_12___mmap_AWQOS),
    .mmap_offset(Mmap2Stream_12___rmem12__q0)
  );


  (* keep_hierarchy = "yes" *) Mmap2Stream
  Mmap2Stream_13
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Mmap2Stream_13__ap_start),
    .ap_done(Mmap2Stream_13__ap_done),
    .ap_idle(Mmap2Stream_13__ap_idle),
    .ap_ready(Mmap2Stream_13__ap_ready),
    .n(Mmap2Stream_13___n__q0),
    .stream_din(qr13_vadd_bw__din),
    .stream_full_n(qr13_vadd_bw__full_n),
    .stream_write(qr13_vadd_bw__write),
    .m_axi_mmap_ARADDR(m_axi_rmem13___Mmap2Stream_13___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem13___Mmap2Stream_13___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem13___Mmap2Stream_13___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem13___Mmap2Stream_13___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem13___Mmap2Stream_13___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem13___Mmap2Stream_13___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem13___Mmap2Stream_13___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem13___Mmap2Stream_13___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem13___Mmap2Stream_13___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem13___Mmap2Stream_13___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem13___Mmap2Stream_13___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem13___Mmap2Stream_13___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem13___Mmap2Stream_13___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem13___Mmap2Stream_13___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem13___Mmap2Stream_13___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem13___Mmap2Stream_13___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem13___Mmap2Stream_13___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem13___Mmap2Stream_13___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem13___Mmap2Stream_13___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem13___Mmap2Stream_13___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem13___Mmap2Stream_13___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem13___Mmap2Stream_13___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem13___Mmap2Stream_13___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem13___Mmap2Stream_13___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem13___Mmap2Stream_13___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem13___Mmap2Stream_13___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem13___Mmap2Stream_13___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem13___Mmap2Stream_13___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem13___Mmap2Stream_13___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem13___Mmap2Stream_13___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem13___Mmap2Stream_13___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem13___Mmap2Stream_13___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem13___Mmap2Stream_13___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem13___Mmap2Stream_13___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem13___Mmap2Stream_13___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem13___Mmap2Stream_13___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem13___Mmap2Stream_13___mmap_AWQOS),
    .mmap_offset(Mmap2Stream_13___rmem13__q0)
  );


  (* keep_hierarchy = "yes" *) Mmap2Stream
  Mmap2Stream_14
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Mmap2Stream_14__ap_start),
    .ap_done(Mmap2Stream_14__ap_done),
    .ap_idle(Mmap2Stream_14__ap_idle),
    .ap_ready(Mmap2Stream_14__ap_ready),
    .n(Mmap2Stream_14___n__q0),
    .stream_din(qr14_vadd_bw__din),
    .stream_full_n(qr14_vadd_bw__full_n),
    .stream_write(qr14_vadd_bw__write),
    .m_axi_mmap_ARADDR(m_axi_rmem14___Mmap2Stream_14___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem14___Mmap2Stream_14___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem14___Mmap2Stream_14___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem14___Mmap2Stream_14___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem14___Mmap2Stream_14___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem14___Mmap2Stream_14___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem14___Mmap2Stream_14___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem14___Mmap2Stream_14___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem14___Mmap2Stream_14___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem14___Mmap2Stream_14___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem14___Mmap2Stream_14___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem14___Mmap2Stream_14___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem14___Mmap2Stream_14___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem14___Mmap2Stream_14___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem14___Mmap2Stream_14___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem14___Mmap2Stream_14___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem14___Mmap2Stream_14___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem14___Mmap2Stream_14___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem14___Mmap2Stream_14___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem14___Mmap2Stream_14___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem14___Mmap2Stream_14___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem14___Mmap2Stream_14___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem14___Mmap2Stream_14___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem14___Mmap2Stream_14___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem14___Mmap2Stream_14___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem14___Mmap2Stream_14___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem14___Mmap2Stream_14___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem14___Mmap2Stream_14___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem14___Mmap2Stream_14___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem14___Mmap2Stream_14___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem14___Mmap2Stream_14___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem14___Mmap2Stream_14___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem14___Mmap2Stream_14___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem14___Mmap2Stream_14___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem14___Mmap2Stream_14___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem14___Mmap2Stream_14___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem14___Mmap2Stream_14___mmap_AWQOS),
    .mmap_offset(Mmap2Stream_14___rmem14__q0)
  );


  (* keep_hierarchy = "yes" *) Mmap2Stream
  Mmap2Stream_15
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Mmap2Stream_15__ap_start),
    .ap_done(Mmap2Stream_15__ap_done),
    .ap_idle(Mmap2Stream_15__ap_idle),
    .ap_ready(Mmap2Stream_15__ap_ready),
    .n(Mmap2Stream_15___n__q0),
    .stream_din(qr15_vadd_bw__din),
    .stream_full_n(qr15_vadd_bw__full_n),
    .stream_write(qr15_vadd_bw__write),
    .m_axi_mmap_ARADDR(m_axi_rmem15___Mmap2Stream_15___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem15___Mmap2Stream_15___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem15___Mmap2Stream_15___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem15___Mmap2Stream_15___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem15___Mmap2Stream_15___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem15___Mmap2Stream_15___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem15___Mmap2Stream_15___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem15___Mmap2Stream_15___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem15___Mmap2Stream_15___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem15___Mmap2Stream_15___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem15___Mmap2Stream_15___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem15___Mmap2Stream_15___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem15___Mmap2Stream_15___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem15___Mmap2Stream_15___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem15___Mmap2Stream_15___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem15___Mmap2Stream_15___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem15___Mmap2Stream_15___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem15___Mmap2Stream_15___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem15___Mmap2Stream_15___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem15___Mmap2Stream_15___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem15___Mmap2Stream_15___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem15___Mmap2Stream_15___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem15___Mmap2Stream_15___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem15___Mmap2Stream_15___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem15___Mmap2Stream_15___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem15___Mmap2Stream_15___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem15___Mmap2Stream_15___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem15___Mmap2Stream_15___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem15___Mmap2Stream_15___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem15___Mmap2Stream_15___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem15___Mmap2Stream_15___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem15___Mmap2Stream_15___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem15___Mmap2Stream_15___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem15___Mmap2Stream_15___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem15___Mmap2Stream_15___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem15___Mmap2Stream_15___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem15___Mmap2Stream_15___mmap_AWQOS),
    .mmap_offset(Mmap2Stream_15___rmem15__q0)
  );


  (* keep_hierarchy = "yes" *) Mmap2Stream
  Mmap2Stream_16
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Mmap2Stream_16__ap_start),
    .ap_done(Mmap2Stream_16__ap_done),
    .ap_idle(Mmap2Stream_16__ap_idle),
    .ap_ready(Mmap2Stream_16__ap_ready),
    .n(Mmap2Stream_16___n__q0),
    .stream_din(qr16_vadd_bw__din),
    .stream_full_n(qr16_vadd_bw__full_n),
    .stream_write(qr16_vadd_bw__write),
    .m_axi_mmap_ARADDR(m_axi_rmem16___Mmap2Stream_16___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem16___Mmap2Stream_16___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem16___Mmap2Stream_16___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem16___Mmap2Stream_16___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem16___Mmap2Stream_16___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem16___Mmap2Stream_16___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem16___Mmap2Stream_16___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem16___Mmap2Stream_16___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem16___Mmap2Stream_16___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem16___Mmap2Stream_16___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem16___Mmap2Stream_16___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem16___Mmap2Stream_16___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem16___Mmap2Stream_16___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem16___Mmap2Stream_16___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem16___Mmap2Stream_16___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem16___Mmap2Stream_16___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem16___Mmap2Stream_16___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem16___Mmap2Stream_16___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem16___Mmap2Stream_16___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem16___Mmap2Stream_16___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem16___Mmap2Stream_16___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem16___Mmap2Stream_16___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem16___Mmap2Stream_16___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem16___Mmap2Stream_16___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem16___Mmap2Stream_16___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem16___Mmap2Stream_16___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem16___Mmap2Stream_16___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem16___Mmap2Stream_16___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem16___Mmap2Stream_16___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem16___Mmap2Stream_16___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem16___Mmap2Stream_16___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem16___Mmap2Stream_16___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem16___Mmap2Stream_16___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem16___Mmap2Stream_16___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem16___Mmap2Stream_16___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem16___Mmap2Stream_16___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem16___Mmap2Stream_16___mmap_AWQOS),
    .mmap_offset(Mmap2Stream_16___rmem16__q0)
  );


  (* keep_hierarchy = "yes" *) Mmap2Stream
  Mmap2Stream_17
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Mmap2Stream_17__ap_start),
    .ap_done(Mmap2Stream_17__ap_done),
    .ap_idle(Mmap2Stream_17__ap_idle),
    .ap_ready(Mmap2Stream_17__ap_ready),
    .n(Mmap2Stream_17___n__q0),
    .stream_din(qr17_vadd_bw__din),
    .stream_full_n(qr17_vadd_bw__full_n),
    .stream_write(qr17_vadd_bw__write),
    .m_axi_mmap_ARADDR(m_axi_rmem17___Mmap2Stream_17___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem17___Mmap2Stream_17___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem17___Mmap2Stream_17___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem17___Mmap2Stream_17___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem17___Mmap2Stream_17___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem17___Mmap2Stream_17___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem17___Mmap2Stream_17___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem17___Mmap2Stream_17___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem17___Mmap2Stream_17___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem17___Mmap2Stream_17___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem17___Mmap2Stream_17___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem17___Mmap2Stream_17___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem17___Mmap2Stream_17___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem17___Mmap2Stream_17___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem17___Mmap2Stream_17___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem17___Mmap2Stream_17___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem17___Mmap2Stream_17___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem17___Mmap2Stream_17___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem17___Mmap2Stream_17___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem17___Mmap2Stream_17___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem17___Mmap2Stream_17___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem17___Mmap2Stream_17___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem17___Mmap2Stream_17___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem17___Mmap2Stream_17___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem17___Mmap2Stream_17___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem17___Mmap2Stream_17___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem17___Mmap2Stream_17___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem17___Mmap2Stream_17___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem17___Mmap2Stream_17___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem17___Mmap2Stream_17___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem17___Mmap2Stream_17___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem17___Mmap2Stream_17___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem17___Mmap2Stream_17___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem17___Mmap2Stream_17___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem17___Mmap2Stream_17___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem17___Mmap2Stream_17___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem17___Mmap2Stream_17___mmap_AWQOS),
    .mmap_offset(Mmap2Stream_17___rmem17__q0)
  );


  (* keep_hierarchy = "yes" *) Mmap2Stream
  Mmap2Stream_18
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Mmap2Stream_18__ap_start),
    .ap_done(Mmap2Stream_18__ap_done),
    .ap_idle(Mmap2Stream_18__ap_idle),
    .ap_ready(Mmap2Stream_18__ap_ready),
    .n(Mmap2Stream_18___n__q0),
    .stream_din(qr18_vadd_bw__din),
    .stream_full_n(qr18_vadd_bw__full_n),
    .stream_write(qr18_vadd_bw__write),
    .m_axi_mmap_ARADDR(m_axi_rmem18___Mmap2Stream_18___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem18___Mmap2Stream_18___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem18___Mmap2Stream_18___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem18___Mmap2Stream_18___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem18___Mmap2Stream_18___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem18___Mmap2Stream_18___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem18___Mmap2Stream_18___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem18___Mmap2Stream_18___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem18___Mmap2Stream_18___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem18___Mmap2Stream_18___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem18___Mmap2Stream_18___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem18___Mmap2Stream_18___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem18___Mmap2Stream_18___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem18___Mmap2Stream_18___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem18___Mmap2Stream_18___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem18___Mmap2Stream_18___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem18___Mmap2Stream_18___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem18___Mmap2Stream_18___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem18___Mmap2Stream_18___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem18___Mmap2Stream_18___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem18___Mmap2Stream_18___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem18___Mmap2Stream_18___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem18___Mmap2Stream_18___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem18___Mmap2Stream_18___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem18___Mmap2Stream_18___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem18___Mmap2Stream_18___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem18___Mmap2Stream_18___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem18___Mmap2Stream_18___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem18___Mmap2Stream_18___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem18___Mmap2Stream_18___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem18___Mmap2Stream_18___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem18___Mmap2Stream_18___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem18___Mmap2Stream_18___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem18___Mmap2Stream_18___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem18___Mmap2Stream_18___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem18___Mmap2Stream_18___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem18___Mmap2Stream_18___mmap_AWQOS),
    .mmap_offset(Mmap2Stream_18___rmem18__q0)
  );


  (* keep_hierarchy = "yes" *) Mmap2Stream
  Mmap2Stream_19
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Mmap2Stream_19__ap_start),
    .ap_done(Mmap2Stream_19__ap_done),
    .ap_idle(Mmap2Stream_19__ap_idle),
    .ap_ready(Mmap2Stream_19__ap_ready),
    .n(Mmap2Stream_19___n__q0),
    .stream_din(qr19_vadd_bw__din),
    .stream_full_n(qr19_vadd_bw__full_n),
    .stream_write(qr19_vadd_bw__write),
    .m_axi_mmap_ARADDR(m_axi_rmem19___Mmap2Stream_19___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem19___Mmap2Stream_19___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem19___Mmap2Stream_19___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem19___Mmap2Stream_19___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem19___Mmap2Stream_19___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem19___Mmap2Stream_19___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem19___Mmap2Stream_19___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem19___Mmap2Stream_19___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem19___Mmap2Stream_19___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem19___Mmap2Stream_19___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem19___Mmap2Stream_19___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem19___Mmap2Stream_19___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem19___Mmap2Stream_19___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem19___Mmap2Stream_19___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem19___Mmap2Stream_19___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem19___Mmap2Stream_19___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem19___Mmap2Stream_19___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem19___Mmap2Stream_19___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem19___Mmap2Stream_19___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem19___Mmap2Stream_19___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem19___Mmap2Stream_19___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem19___Mmap2Stream_19___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem19___Mmap2Stream_19___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem19___Mmap2Stream_19___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem19___Mmap2Stream_19___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem19___Mmap2Stream_19___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem19___Mmap2Stream_19___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem19___Mmap2Stream_19___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem19___Mmap2Stream_19___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem19___Mmap2Stream_19___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem19___Mmap2Stream_19___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem19___Mmap2Stream_19___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem19___Mmap2Stream_19___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem19___Mmap2Stream_19___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem19___Mmap2Stream_19___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem19___Mmap2Stream_19___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem19___Mmap2Stream_19___mmap_AWQOS),
    .mmap_offset(Mmap2Stream_19___rmem19__q0)
  );


  (* keep_hierarchy = "yes" *) Mmap2Stream
  Mmap2Stream_20
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Mmap2Stream_20__ap_start),
    .ap_done(Mmap2Stream_20__ap_done),
    .ap_idle(Mmap2Stream_20__ap_idle),
    .ap_ready(Mmap2Stream_20__ap_ready),
    .n(Mmap2Stream_20___n__q0),
    .stream_din(qr20_vadd_bw__din),
    .stream_full_n(qr20_vadd_bw__full_n),
    .stream_write(qr20_vadd_bw__write),
    .m_axi_mmap_ARADDR(m_axi_rmem20___Mmap2Stream_20___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem20___Mmap2Stream_20___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem20___Mmap2Stream_20___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem20___Mmap2Stream_20___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem20___Mmap2Stream_20___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem20___Mmap2Stream_20___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem20___Mmap2Stream_20___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem20___Mmap2Stream_20___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem20___Mmap2Stream_20___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem20___Mmap2Stream_20___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem20___Mmap2Stream_20___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem20___Mmap2Stream_20___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem20___Mmap2Stream_20___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem20___Mmap2Stream_20___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem20___Mmap2Stream_20___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem20___Mmap2Stream_20___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem20___Mmap2Stream_20___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem20___Mmap2Stream_20___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem20___Mmap2Stream_20___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem20___Mmap2Stream_20___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem20___Mmap2Stream_20___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem20___Mmap2Stream_20___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem20___Mmap2Stream_20___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem20___Mmap2Stream_20___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem20___Mmap2Stream_20___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem20___Mmap2Stream_20___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem20___Mmap2Stream_20___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem20___Mmap2Stream_20___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem20___Mmap2Stream_20___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem20___Mmap2Stream_20___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem20___Mmap2Stream_20___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem20___Mmap2Stream_20___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem20___Mmap2Stream_20___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem20___Mmap2Stream_20___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem20___Mmap2Stream_20___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem20___Mmap2Stream_20___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem20___Mmap2Stream_20___mmap_AWQOS),
    .mmap_offset(Mmap2Stream_20___rmem20__q0)
  );


  (* keep_hierarchy = "yes" *) Mmap2Stream
  Mmap2Stream_21
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Mmap2Stream_21__ap_start),
    .ap_done(Mmap2Stream_21__ap_done),
    .ap_idle(Mmap2Stream_21__ap_idle),
    .ap_ready(Mmap2Stream_21__ap_ready),
    .n(Mmap2Stream_21___n__q0),
    .stream_din(qr21_vadd_bw__din),
    .stream_full_n(qr21_vadd_bw__full_n),
    .stream_write(qr21_vadd_bw__write),
    .m_axi_mmap_ARADDR(m_axi_rmem21___Mmap2Stream_21___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem21___Mmap2Stream_21___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem21___Mmap2Stream_21___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem21___Mmap2Stream_21___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem21___Mmap2Stream_21___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem21___Mmap2Stream_21___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem21___Mmap2Stream_21___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem21___Mmap2Stream_21___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem21___Mmap2Stream_21___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem21___Mmap2Stream_21___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem21___Mmap2Stream_21___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem21___Mmap2Stream_21___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem21___Mmap2Stream_21___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem21___Mmap2Stream_21___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem21___Mmap2Stream_21___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem21___Mmap2Stream_21___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem21___Mmap2Stream_21___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem21___Mmap2Stream_21___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem21___Mmap2Stream_21___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem21___Mmap2Stream_21___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem21___Mmap2Stream_21___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem21___Mmap2Stream_21___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem21___Mmap2Stream_21___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem21___Mmap2Stream_21___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem21___Mmap2Stream_21___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem21___Mmap2Stream_21___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem21___Mmap2Stream_21___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem21___Mmap2Stream_21___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem21___Mmap2Stream_21___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem21___Mmap2Stream_21___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem21___Mmap2Stream_21___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem21___Mmap2Stream_21___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem21___Mmap2Stream_21___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem21___Mmap2Stream_21___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem21___Mmap2Stream_21___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem21___Mmap2Stream_21___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem21___Mmap2Stream_21___mmap_AWQOS),
    .mmap_offset(Mmap2Stream_21___rmem21__q0)
  );


  (* keep_hierarchy = "yes" *) Mmap2Stream
  Mmap2Stream_22
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Mmap2Stream_22__ap_start),
    .ap_done(Mmap2Stream_22__ap_done),
    .ap_idle(Mmap2Stream_22__ap_idle),
    .ap_ready(Mmap2Stream_22__ap_ready),
    .n(Mmap2Stream_22___n__q0),
    .stream_din(qr22_vadd_bw__din),
    .stream_full_n(qr22_vadd_bw__full_n),
    .stream_write(qr22_vadd_bw__write),
    .m_axi_mmap_ARADDR(m_axi_rmem22___Mmap2Stream_22___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem22___Mmap2Stream_22___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem22___Mmap2Stream_22___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem22___Mmap2Stream_22___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem22___Mmap2Stream_22___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem22___Mmap2Stream_22___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem22___Mmap2Stream_22___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem22___Mmap2Stream_22___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem22___Mmap2Stream_22___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem22___Mmap2Stream_22___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem22___Mmap2Stream_22___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem22___Mmap2Stream_22___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem22___Mmap2Stream_22___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem22___Mmap2Stream_22___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem22___Mmap2Stream_22___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem22___Mmap2Stream_22___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem22___Mmap2Stream_22___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem22___Mmap2Stream_22___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem22___Mmap2Stream_22___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem22___Mmap2Stream_22___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem22___Mmap2Stream_22___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem22___Mmap2Stream_22___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem22___Mmap2Stream_22___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem22___Mmap2Stream_22___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem22___Mmap2Stream_22___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem22___Mmap2Stream_22___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem22___Mmap2Stream_22___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem22___Mmap2Stream_22___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem22___Mmap2Stream_22___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem22___Mmap2Stream_22___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem22___Mmap2Stream_22___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem22___Mmap2Stream_22___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem22___Mmap2Stream_22___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem22___Mmap2Stream_22___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem22___Mmap2Stream_22___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem22___Mmap2Stream_22___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem22___Mmap2Stream_22___mmap_AWQOS),
    .mmap_offset(Mmap2Stream_22___rmem22__q0)
  );


  (* keep_hierarchy = "yes" *) Mmap2Stream
  Mmap2Stream_23
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Mmap2Stream_23__ap_start),
    .ap_done(Mmap2Stream_23__ap_done),
    .ap_idle(Mmap2Stream_23__ap_idle),
    .ap_ready(Mmap2Stream_23__ap_ready),
    .n(Mmap2Stream_23___n__q0),
    .stream_din(qr23_vadd_bw__din),
    .stream_full_n(qr23_vadd_bw__full_n),
    .stream_write(qr23_vadd_bw__write),
    .m_axi_mmap_ARADDR(m_axi_rmem23___Mmap2Stream_23___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem23___Mmap2Stream_23___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem23___Mmap2Stream_23___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem23___Mmap2Stream_23___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem23___Mmap2Stream_23___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem23___Mmap2Stream_23___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem23___Mmap2Stream_23___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem23___Mmap2Stream_23___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem23___Mmap2Stream_23___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem23___Mmap2Stream_23___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem23___Mmap2Stream_23___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem23___Mmap2Stream_23___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem23___Mmap2Stream_23___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem23___Mmap2Stream_23___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem23___Mmap2Stream_23___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem23___Mmap2Stream_23___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem23___Mmap2Stream_23___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem23___Mmap2Stream_23___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem23___Mmap2Stream_23___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem23___Mmap2Stream_23___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem23___Mmap2Stream_23___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem23___Mmap2Stream_23___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem23___Mmap2Stream_23___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem23___Mmap2Stream_23___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem23___Mmap2Stream_23___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem23___Mmap2Stream_23___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem23___Mmap2Stream_23___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem23___Mmap2Stream_23___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem23___Mmap2Stream_23___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem23___Mmap2Stream_23___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem23___Mmap2Stream_23___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem23___Mmap2Stream_23___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem23___Mmap2Stream_23___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem23___Mmap2Stream_23___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem23___Mmap2Stream_23___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem23___Mmap2Stream_23___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem23___Mmap2Stream_23___mmap_AWQOS),
    .mmap_offset(Mmap2Stream_23___rmem23__q0)
  );


  (* keep_hierarchy = "yes" *) Mmap2Stream
  Mmap2Stream_24
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Mmap2Stream_24__ap_start),
    .ap_done(Mmap2Stream_24__ap_done),
    .ap_idle(Mmap2Stream_24__ap_idle),
    .ap_ready(Mmap2Stream_24__ap_ready),
    .n(Mmap2Stream_24___n__q0),
    .stream_din(qr24_vadd_bw__din),
    .stream_full_n(qr24_vadd_bw__full_n),
    .stream_write(qr24_vadd_bw__write),
    .m_axi_mmap_ARADDR(m_axi_rmem24___Mmap2Stream_24___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem24___Mmap2Stream_24___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem24___Mmap2Stream_24___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem24___Mmap2Stream_24___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem24___Mmap2Stream_24___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem24___Mmap2Stream_24___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem24___Mmap2Stream_24___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem24___Mmap2Stream_24___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem24___Mmap2Stream_24___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem24___Mmap2Stream_24___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem24___Mmap2Stream_24___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem24___Mmap2Stream_24___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem24___Mmap2Stream_24___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem24___Mmap2Stream_24___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem24___Mmap2Stream_24___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem24___Mmap2Stream_24___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem24___Mmap2Stream_24___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem24___Mmap2Stream_24___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem24___Mmap2Stream_24___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem24___Mmap2Stream_24___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem24___Mmap2Stream_24___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem24___Mmap2Stream_24___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem24___Mmap2Stream_24___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem24___Mmap2Stream_24___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem24___Mmap2Stream_24___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem24___Mmap2Stream_24___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem24___Mmap2Stream_24___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem24___Mmap2Stream_24___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem24___Mmap2Stream_24___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem24___Mmap2Stream_24___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem24___Mmap2Stream_24___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem24___Mmap2Stream_24___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem24___Mmap2Stream_24___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem24___Mmap2Stream_24___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem24___Mmap2Stream_24___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem24___Mmap2Stream_24___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem24___Mmap2Stream_24___mmap_AWQOS),
    .mmap_offset(Mmap2Stream_24___rmem24__q0)
  );


  (* keep_hierarchy = "yes" *) Mmap2Stream
  Mmap2Stream_25
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Mmap2Stream_25__ap_start),
    .ap_done(Mmap2Stream_25__ap_done),
    .ap_idle(Mmap2Stream_25__ap_idle),
    .ap_ready(Mmap2Stream_25__ap_ready),
    .n(Mmap2Stream_25___n__q0),
    .stream_din(qr25_vadd_bw__din),
    .stream_full_n(qr25_vadd_bw__full_n),
    .stream_write(qr25_vadd_bw__write),
    .m_axi_mmap_ARADDR(m_axi_rmem25___Mmap2Stream_25___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem25___Mmap2Stream_25___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem25___Mmap2Stream_25___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem25___Mmap2Stream_25___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem25___Mmap2Stream_25___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem25___Mmap2Stream_25___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem25___Mmap2Stream_25___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem25___Mmap2Stream_25___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem25___Mmap2Stream_25___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem25___Mmap2Stream_25___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem25___Mmap2Stream_25___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem25___Mmap2Stream_25___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem25___Mmap2Stream_25___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem25___Mmap2Stream_25___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem25___Mmap2Stream_25___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem25___Mmap2Stream_25___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem25___Mmap2Stream_25___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem25___Mmap2Stream_25___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem25___Mmap2Stream_25___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem25___Mmap2Stream_25___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem25___Mmap2Stream_25___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem25___Mmap2Stream_25___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem25___Mmap2Stream_25___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem25___Mmap2Stream_25___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem25___Mmap2Stream_25___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem25___Mmap2Stream_25___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem25___Mmap2Stream_25___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem25___Mmap2Stream_25___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem25___Mmap2Stream_25___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem25___Mmap2Stream_25___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem25___Mmap2Stream_25___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem25___Mmap2Stream_25___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem25___Mmap2Stream_25___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem25___Mmap2Stream_25___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem25___Mmap2Stream_25___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem25___Mmap2Stream_25___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem25___Mmap2Stream_25___mmap_AWQOS),
    .mmap_offset(Mmap2Stream_25___rmem25__q0)
  );


  (* keep_hierarchy = "yes" *) Mmap2Stream
  Mmap2Stream_26
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Mmap2Stream_26__ap_start),
    .ap_done(Mmap2Stream_26__ap_done),
    .ap_idle(Mmap2Stream_26__ap_idle),
    .ap_ready(Mmap2Stream_26__ap_ready),
    .n(Mmap2Stream_26___n__q0),
    .stream_din(qr26_vadd_bw__din),
    .stream_full_n(qr26_vadd_bw__full_n),
    .stream_write(qr26_vadd_bw__write),
    .m_axi_mmap_ARADDR(m_axi_rmem26___Mmap2Stream_26___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem26___Mmap2Stream_26___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem26___Mmap2Stream_26___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem26___Mmap2Stream_26___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem26___Mmap2Stream_26___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem26___Mmap2Stream_26___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem26___Mmap2Stream_26___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem26___Mmap2Stream_26___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem26___Mmap2Stream_26___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem26___Mmap2Stream_26___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem26___Mmap2Stream_26___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem26___Mmap2Stream_26___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem26___Mmap2Stream_26___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem26___Mmap2Stream_26___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem26___Mmap2Stream_26___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem26___Mmap2Stream_26___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem26___Mmap2Stream_26___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem26___Mmap2Stream_26___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem26___Mmap2Stream_26___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem26___Mmap2Stream_26___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem26___Mmap2Stream_26___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem26___Mmap2Stream_26___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem26___Mmap2Stream_26___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem26___Mmap2Stream_26___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem26___Mmap2Stream_26___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem26___Mmap2Stream_26___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem26___Mmap2Stream_26___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem26___Mmap2Stream_26___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem26___Mmap2Stream_26___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem26___Mmap2Stream_26___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem26___Mmap2Stream_26___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem26___Mmap2Stream_26___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem26___Mmap2Stream_26___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem26___Mmap2Stream_26___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem26___Mmap2Stream_26___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem26___Mmap2Stream_26___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem26___Mmap2Stream_26___mmap_AWQOS),
    .mmap_offset(Mmap2Stream_26___rmem26__q0)
  );


  (* keep_hierarchy = "yes" *) Mmap2Stream
  Mmap2Stream_27
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Mmap2Stream_27__ap_start),
    .ap_done(Mmap2Stream_27__ap_done),
    .ap_idle(Mmap2Stream_27__ap_idle),
    .ap_ready(Mmap2Stream_27__ap_ready),
    .n(Mmap2Stream_27___n__q0),
    .stream_din(qr27_vadd_bw__din),
    .stream_full_n(qr27_vadd_bw__full_n),
    .stream_write(qr27_vadd_bw__write),
    .m_axi_mmap_ARADDR(m_axi_rmem27___Mmap2Stream_27___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem27___Mmap2Stream_27___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem27___Mmap2Stream_27___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem27___Mmap2Stream_27___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem27___Mmap2Stream_27___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem27___Mmap2Stream_27___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem27___Mmap2Stream_27___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem27___Mmap2Stream_27___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem27___Mmap2Stream_27___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem27___Mmap2Stream_27___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem27___Mmap2Stream_27___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem27___Mmap2Stream_27___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem27___Mmap2Stream_27___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem27___Mmap2Stream_27___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem27___Mmap2Stream_27___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem27___Mmap2Stream_27___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem27___Mmap2Stream_27___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem27___Mmap2Stream_27___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem27___Mmap2Stream_27___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem27___Mmap2Stream_27___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem27___Mmap2Stream_27___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem27___Mmap2Stream_27___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem27___Mmap2Stream_27___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem27___Mmap2Stream_27___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem27___Mmap2Stream_27___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem27___Mmap2Stream_27___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem27___Mmap2Stream_27___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem27___Mmap2Stream_27___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem27___Mmap2Stream_27___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem27___Mmap2Stream_27___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem27___Mmap2Stream_27___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem27___Mmap2Stream_27___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem27___Mmap2Stream_27___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem27___Mmap2Stream_27___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem27___Mmap2Stream_27___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem27___Mmap2Stream_27___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem27___Mmap2Stream_27___mmap_AWQOS),
    .mmap_offset(Mmap2Stream_27___rmem27__q0)
  );


  (* keep_hierarchy = "yes" *) Stream2Mmap
  Stream2Mmap_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Stream2Mmap_0__ap_start),
    .ap_done(Stream2Mmap_0__ap_done),
    .ap_idle(Stream2Mmap_0__ap_idle),
    .ap_ready(Stream2Mmap_0__ap_ready),
    .n(Stream2Mmap_0___n__q0),
    .stream_s_dout(qw0_vadd_bw__dout),
    .stream_peek_dout(qw0_vadd_bw__dout),
    .stream_s_empty_n(qw0_vadd_bw__empty_n),
    .stream_peek_empty_n(qw0_vadd_bw__empty_n),
    .stream_s_read(qw0_vadd_bw__read),
    .stream_peek_read(),
    .m_axi_mmap_ARADDR(m_axi_rmem0___Stream2Mmap_0___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem0___Stream2Mmap_0___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem0___Stream2Mmap_0___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem0___Stream2Mmap_0___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem0___Stream2Mmap_0___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem0___Stream2Mmap_0___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem0___Stream2Mmap_0___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem0___Stream2Mmap_0___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem0___Stream2Mmap_0___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem0___Stream2Mmap_0___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem0___Stream2Mmap_0___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem0___Stream2Mmap_0___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem0___Stream2Mmap_0___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem0___Stream2Mmap_0___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem0___Stream2Mmap_0___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem0___Stream2Mmap_0___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem0___Stream2Mmap_0___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem0___Stream2Mmap_0___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem0___Stream2Mmap_0___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem0___Stream2Mmap_0___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem0___Stream2Mmap_0___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem0___Stream2Mmap_0___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem0___Stream2Mmap_0___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem0___Stream2Mmap_0___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem0___Stream2Mmap_0___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem0___Stream2Mmap_0___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem0___Stream2Mmap_0___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem0___Stream2Mmap_0___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem0___Stream2Mmap_0___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem0___Stream2Mmap_0___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem0___Stream2Mmap_0___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem0___Stream2Mmap_0___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem0___Stream2Mmap_0___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem0___Stream2Mmap_0___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem0___Stream2Mmap_0___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem0___Stream2Mmap_0___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem0___Stream2Mmap_0___mmap_AWQOS),
    .mmap_offset(Stream2Mmap_0___rmem0__q0)
  );


  (* keep_hierarchy = "yes" *) Stream2Mmap
  Stream2Mmap_1
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Stream2Mmap_1__ap_start),
    .ap_done(Stream2Mmap_1__ap_done),
    .ap_idle(Stream2Mmap_1__ap_idle),
    .ap_ready(Stream2Mmap_1__ap_ready),
    .n(Stream2Mmap_1___n__q0),
    .stream_s_dout(qw1_vadd_bw__dout),
    .stream_peek_dout(qw1_vadd_bw__dout),
    .stream_s_empty_n(qw1_vadd_bw__empty_n),
    .stream_peek_empty_n(qw1_vadd_bw__empty_n),
    .stream_s_read(qw1_vadd_bw__read),
    .stream_peek_read(),
    .m_axi_mmap_ARADDR(m_axi_rmem1___Stream2Mmap_1___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem1___Stream2Mmap_1___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem1___Stream2Mmap_1___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem1___Stream2Mmap_1___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem1___Stream2Mmap_1___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem1___Stream2Mmap_1___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem1___Stream2Mmap_1___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem1___Stream2Mmap_1___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem1___Stream2Mmap_1___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem1___Stream2Mmap_1___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem1___Stream2Mmap_1___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem1___Stream2Mmap_1___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem1___Stream2Mmap_1___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem1___Stream2Mmap_1___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem1___Stream2Mmap_1___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem1___Stream2Mmap_1___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem1___Stream2Mmap_1___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem1___Stream2Mmap_1___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem1___Stream2Mmap_1___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem1___Stream2Mmap_1___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem1___Stream2Mmap_1___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem1___Stream2Mmap_1___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem1___Stream2Mmap_1___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem1___Stream2Mmap_1___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem1___Stream2Mmap_1___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem1___Stream2Mmap_1___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem1___Stream2Mmap_1___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem1___Stream2Mmap_1___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem1___Stream2Mmap_1___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem1___Stream2Mmap_1___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem1___Stream2Mmap_1___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem1___Stream2Mmap_1___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem1___Stream2Mmap_1___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem1___Stream2Mmap_1___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem1___Stream2Mmap_1___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem1___Stream2Mmap_1___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem1___Stream2Mmap_1___mmap_AWQOS),
    .mmap_offset(Stream2Mmap_1___rmem1__q0)
  );


  (* keep_hierarchy = "yes" *) Stream2Mmap
  Stream2Mmap_2
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Stream2Mmap_2__ap_start),
    .ap_done(Stream2Mmap_2__ap_done),
    .ap_idle(Stream2Mmap_2__ap_idle),
    .ap_ready(Stream2Mmap_2__ap_ready),
    .n(Stream2Mmap_2___n__q0),
    .stream_s_dout(qw2_vadd_bw__dout),
    .stream_peek_dout(qw2_vadd_bw__dout),
    .stream_s_empty_n(qw2_vadd_bw__empty_n),
    .stream_peek_empty_n(qw2_vadd_bw__empty_n),
    .stream_s_read(qw2_vadd_bw__read),
    .stream_peek_read(),
    .m_axi_mmap_ARADDR(m_axi_rmem2___Stream2Mmap_2___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem2___Stream2Mmap_2___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem2___Stream2Mmap_2___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem2___Stream2Mmap_2___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem2___Stream2Mmap_2___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem2___Stream2Mmap_2___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem2___Stream2Mmap_2___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem2___Stream2Mmap_2___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem2___Stream2Mmap_2___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem2___Stream2Mmap_2___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem2___Stream2Mmap_2___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem2___Stream2Mmap_2___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem2___Stream2Mmap_2___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem2___Stream2Mmap_2___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem2___Stream2Mmap_2___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem2___Stream2Mmap_2___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem2___Stream2Mmap_2___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem2___Stream2Mmap_2___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem2___Stream2Mmap_2___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem2___Stream2Mmap_2___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem2___Stream2Mmap_2___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem2___Stream2Mmap_2___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem2___Stream2Mmap_2___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem2___Stream2Mmap_2___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem2___Stream2Mmap_2___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem2___Stream2Mmap_2___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem2___Stream2Mmap_2___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem2___Stream2Mmap_2___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem2___Stream2Mmap_2___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem2___Stream2Mmap_2___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem2___Stream2Mmap_2___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem2___Stream2Mmap_2___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem2___Stream2Mmap_2___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem2___Stream2Mmap_2___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem2___Stream2Mmap_2___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem2___Stream2Mmap_2___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem2___Stream2Mmap_2___mmap_AWQOS),
    .mmap_offset(Stream2Mmap_2___rmem2__q0)
  );


  (* keep_hierarchy = "yes" *) Stream2Mmap
  Stream2Mmap_3
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Stream2Mmap_3__ap_start),
    .ap_done(Stream2Mmap_3__ap_done),
    .ap_idle(Stream2Mmap_3__ap_idle),
    .ap_ready(Stream2Mmap_3__ap_ready),
    .n(Stream2Mmap_3___n__q0),
    .stream_s_dout(qw3_vadd_bw__dout),
    .stream_peek_dout(qw3_vadd_bw__dout),
    .stream_s_empty_n(qw3_vadd_bw__empty_n),
    .stream_peek_empty_n(qw3_vadd_bw__empty_n),
    .stream_s_read(qw3_vadd_bw__read),
    .stream_peek_read(),
    .m_axi_mmap_ARADDR(m_axi_rmem3___Stream2Mmap_3___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem3___Stream2Mmap_3___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem3___Stream2Mmap_3___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem3___Stream2Mmap_3___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem3___Stream2Mmap_3___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem3___Stream2Mmap_3___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem3___Stream2Mmap_3___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem3___Stream2Mmap_3___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem3___Stream2Mmap_3___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem3___Stream2Mmap_3___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem3___Stream2Mmap_3___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem3___Stream2Mmap_3___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem3___Stream2Mmap_3___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem3___Stream2Mmap_3___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem3___Stream2Mmap_3___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem3___Stream2Mmap_3___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem3___Stream2Mmap_3___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem3___Stream2Mmap_3___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem3___Stream2Mmap_3___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem3___Stream2Mmap_3___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem3___Stream2Mmap_3___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem3___Stream2Mmap_3___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem3___Stream2Mmap_3___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem3___Stream2Mmap_3___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem3___Stream2Mmap_3___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem3___Stream2Mmap_3___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem3___Stream2Mmap_3___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem3___Stream2Mmap_3___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem3___Stream2Mmap_3___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem3___Stream2Mmap_3___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem3___Stream2Mmap_3___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem3___Stream2Mmap_3___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem3___Stream2Mmap_3___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem3___Stream2Mmap_3___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem3___Stream2Mmap_3___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem3___Stream2Mmap_3___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem3___Stream2Mmap_3___mmap_AWQOS),
    .mmap_offset(Stream2Mmap_3___rmem3__q0)
  );


  (* keep_hierarchy = "yes" *) Stream2Mmap
  Stream2Mmap_4
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Stream2Mmap_4__ap_start),
    .ap_done(Stream2Mmap_4__ap_done),
    .ap_idle(Stream2Mmap_4__ap_idle),
    .ap_ready(Stream2Mmap_4__ap_ready),
    .n(Stream2Mmap_4___n__q0),
    .stream_s_dout(qw4_vadd_bw__dout),
    .stream_peek_dout(qw4_vadd_bw__dout),
    .stream_s_empty_n(qw4_vadd_bw__empty_n),
    .stream_peek_empty_n(qw4_vadd_bw__empty_n),
    .stream_s_read(qw4_vadd_bw__read),
    .stream_peek_read(),
    .m_axi_mmap_ARADDR(m_axi_rmem4___Stream2Mmap_4___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem4___Stream2Mmap_4___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem4___Stream2Mmap_4___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem4___Stream2Mmap_4___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem4___Stream2Mmap_4___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem4___Stream2Mmap_4___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem4___Stream2Mmap_4___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem4___Stream2Mmap_4___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem4___Stream2Mmap_4___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem4___Stream2Mmap_4___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem4___Stream2Mmap_4___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem4___Stream2Mmap_4___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem4___Stream2Mmap_4___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem4___Stream2Mmap_4___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem4___Stream2Mmap_4___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem4___Stream2Mmap_4___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem4___Stream2Mmap_4___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem4___Stream2Mmap_4___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem4___Stream2Mmap_4___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem4___Stream2Mmap_4___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem4___Stream2Mmap_4___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem4___Stream2Mmap_4___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem4___Stream2Mmap_4___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem4___Stream2Mmap_4___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem4___Stream2Mmap_4___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem4___Stream2Mmap_4___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem4___Stream2Mmap_4___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem4___Stream2Mmap_4___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem4___Stream2Mmap_4___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem4___Stream2Mmap_4___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem4___Stream2Mmap_4___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem4___Stream2Mmap_4___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem4___Stream2Mmap_4___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem4___Stream2Mmap_4___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem4___Stream2Mmap_4___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem4___Stream2Mmap_4___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem4___Stream2Mmap_4___mmap_AWQOS),
    .mmap_offset(Stream2Mmap_4___rmem4__q0)
  );


  (* keep_hierarchy = "yes" *) Stream2Mmap
  Stream2Mmap_5
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Stream2Mmap_5__ap_start),
    .ap_done(Stream2Mmap_5__ap_done),
    .ap_idle(Stream2Mmap_5__ap_idle),
    .ap_ready(Stream2Mmap_5__ap_ready),
    .n(Stream2Mmap_5___n__q0),
    .stream_s_dout(qw5_vadd_bw__dout),
    .stream_peek_dout(qw5_vadd_bw__dout),
    .stream_s_empty_n(qw5_vadd_bw__empty_n),
    .stream_peek_empty_n(qw5_vadd_bw__empty_n),
    .stream_s_read(qw5_vadd_bw__read),
    .stream_peek_read(),
    .m_axi_mmap_ARADDR(m_axi_rmem5___Stream2Mmap_5___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem5___Stream2Mmap_5___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem5___Stream2Mmap_5___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem5___Stream2Mmap_5___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem5___Stream2Mmap_5___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem5___Stream2Mmap_5___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem5___Stream2Mmap_5___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem5___Stream2Mmap_5___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem5___Stream2Mmap_5___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem5___Stream2Mmap_5___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem5___Stream2Mmap_5___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem5___Stream2Mmap_5___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem5___Stream2Mmap_5___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem5___Stream2Mmap_5___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem5___Stream2Mmap_5___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem5___Stream2Mmap_5___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem5___Stream2Mmap_5___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem5___Stream2Mmap_5___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem5___Stream2Mmap_5___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem5___Stream2Mmap_5___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem5___Stream2Mmap_5___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem5___Stream2Mmap_5___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem5___Stream2Mmap_5___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem5___Stream2Mmap_5___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem5___Stream2Mmap_5___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem5___Stream2Mmap_5___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem5___Stream2Mmap_5___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem5___Stream2Mmap_5___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem5___Stream2Mmap_5___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem5___Stream2Mmap_5___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem5___Stream2Mmap_5___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem5___Stream2Mmap_5___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem5___Stream2Mmap_5___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem5___Stream2Mmap_5___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem5___Stream2Mmap_5___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem5___Stream2Mmap_5___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem5___Stream2Mmap_5___mmap_AWQOS),
    .mmap_offset(Stream2Mmap_5___rmem5__q0)
  );


  (* keep_hierarchy = "yes" *) Stream2Mmap
  Stream2Mmap_6
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Stream2Mmap_6__ap_start),
    .ap_done(Stream2Mmap_6__ap_done),
    .ap_idle(Stream2Mmap_6__ap_idle),
    .ap_ready(Stream2Mmap_6__ap_ready),
    .n(Stream2Mmap_6___n__q0),
    .stream_s_dout(qw6_vadd_bw__dout),
    .stream_peek_dout(qw6_vadd_bw__dout),
    .stream_s_empty_n(qw6_vadd_bw__empty_n),
    .stream_peek_empty_n(qw6_vadd_bw__empty_n),
    .stream_s_read(qw6_vadd_bw__read),
    .stream_peek_read(),
    .m_axi_mmap_ARADDR(m_axi_rmem6___Stream2Mmap_6___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem6___Stream2Mmap_6___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem6___Stream2Mmap_6___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem6___Stream2Mmap_6___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem6___Stream2Mmap_6___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem6___Stream2Mmap_6___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem6___Stream2Mmap_6___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem6___Stream2Mmap_6___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem6___Stream2Mmap_6___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem6___Stream2Mmap_6___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem6___Stream2Mmap_6___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem6___Stream2Mmap_6___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem6___Stream2Mmap_6___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem6___Stream2Mmap_6___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem6___Stream2Mmap_6___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem6___Stream2Mmap_6___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem6___Stream2Mmap_6___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem6___Stream2Mmap_6___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem6___Stream2Mmap_6___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem6___Stream2Mmap_6___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem6___Stream2Mmap_6___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem6___Stream2Mmap_6___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem6___Stream2Mmap_6___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem6___Stream2Mmap_6___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem6___Stream2Mmap_6___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem6___Stream2Mmap_6___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem6___Stream2Mmap_6___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem6___Stream2Mmap_6___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem6___Stream2Mmap_6___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem6___Stream2Mmap_6___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem6___Stream2Mmap_6___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem6___Stream2Mmap_6___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem6___Stream2Mmap_6___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem6___Stream2Mmap_6___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem6___Stream2Mmap_6___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem6___Stream2Mmap_6___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem6___Stream2Mmap_6___mmap_AWQOS),
    .mmap_offset(Stream2Mmap_6___rmem6__q0)
  );


  (* keep_hierarchy = "yes" *) Stream2Mmap
  Stream2Mmap_7
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Stream2Mmap_7__ap_start),
    .ap_done(Stream2Mmap_7__ap_done),
    .ap_idle(Stream2Mmap_7__ap_idle),
    .ap_ready(Stream2Mmap_7__ap_ready),
    .n(Stream2Mmap_7___n__q0),
    .stream_s_dout(qw7_vadd_bw__dout),
    .stream_peek_dout(qw7_vadd_bw__dout),
    .stream_s_empty_n(qw7_vadd_bw__empty_n),
    .stream_peek_empty_n(qw7_vadd_bw__empty_n),
    .stream_s_read(qw7_vadd_bw__read),
    .stream_peek_read(),
    .m_axi_mmap_ARADDR(m_axi_rmem7___Stream2Mmap_7___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem7___Stream2Mmap_7___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem7___Stream2Mmap_7___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem7___Stream2Mmap_7___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem7___Stream2Mmap_7___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem7___Stream2Mmap_7___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem7___Stream2Mmap_7___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem7___Stream2Mmap_7___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem7___Stream2Mmap_7___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem7___Stream2Mmap_7___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem7___Stream2Mmap_7___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem7___Stream2Mmap_7___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem7___Stream2Mmap_7___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem7___Stream2Mmap_7___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem7___Stream2Mmap_7___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem7___Stream2Mmap_7___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem7___Stream2Mmap_7___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem7___Stream2Mmap_7___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem7___Stream2Mmap_7___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem7___Stream2Mmap_7___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem7___Stream2Mmap_7___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem7___Stream2Mmap_7___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem7___Stream2Mmap_7___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem7___Stream2Mmap_7___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem7___Stream2Mmap_7___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem7___Stream2Mmap_7___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem7___Stream2Mmap_7___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem7___Stream2Mmap_7___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem7___Stream2Mmap_7___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem7___Stream2Mmap_7___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem7___Stream2Mmap_7___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem7___Stream2Mmap_7___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem7___Stream2Mmap_7___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem7___Stream2Mmap_7___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem7___Stream2Mmap_7___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem7___Stream2Mmap_7___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem7___Stream2Mmap_7___mmap_AWQOS),
    .mmap_offset(Stream2Mmap_7___rmem7__q0)
  );


  (* keep_hierarchy = "yes" *) Stream2Mmap
  Stream2Mmap_8
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Stream2Mmap_8__ap_start),
    .ap_done(Stream2Mmap_8__ap_done),
    .ap_idle(Stream2Mmap_8__ap_idle),
    .ap_ready(Stream2Mmap_8__ap_ready),
    .n(Stream2Mmap_8___n__q0),
    .stream_s_dout(qw8_vadd_bw__dout),
    .stream_peek_dout(qw8_vadd_bw__dout),
    .stream_s_empty_n(qw8_vadd_bw__empty_n),
    .stream_peek_empty_n(qw8_vadd_bw__empty_n),
    .stream_s_read(qw8_vadd_bw__read),
    .stream_peek_read(),
    .m_axi_mmap_ARADDR(m_axi_rmem8___Stream2Mmap_8___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem8___Stream2Mmap_8___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem8___Stream2Mmap_8___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem8___Stream2Mmap_8___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem8___Stream2Mmap_8___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem8___Stream2Mmap_8___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem8___Stream2Mmap_8___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem8___Stream2Mmap_8___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem8___Stream2Mmap_8___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem8___Stream2Mmap_8___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem8___Stream2Mmap_8___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem8___Stream2Mmap_8___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem8___Stream2Mmap_8___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem8___Stream2Mmap_8___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem8___Stream2Mmap_8___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem8___Stream2Mmap_8___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem8___Stream2Mmap_8___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem8___Stream2Mmap_8___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem8___Stream2Mmap_8___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem8___Stream2Mmap_8___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem8___Stream2Mmap_8___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem8___Stream2Mmap_8___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem8___Stream2Mmap_8___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem8___Stream2Mmap_8___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem8___Stream2Mmap_8___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem8___Stream2Mmap_8___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem8___Stream2Mmap_8___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem8___Stream2Mmap_8___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem8___Stream2Mmap_8___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem8___Stream2Mmap_8___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem8___Stream2Mmap_8___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem8___Stream2Mmap_8___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem8___Stream2Mmap_8___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem8___Stream2Mmap_8___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem8___Stream2Mmap_8___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem8___Stream2Mmap_8___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem8___Stream2Mmap_8___mmap_AWQOS),
    .mmap_offset(Stream2Mmap_8___rmem8__q0)
  );


  (* keep_hierarchy = "yes" *) Stream2Mmap
  Stream2Mmap_9
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Stream2Mmap_9__ap_start),
    .ap_done(Stream2Mmap_9__ap_done),
    .ap_idle(Stream2Mmap_9__ap_idle),
    .ap_ready(Stream2Mmap_9__ap_ready),
    .n(Stream2Mmap_9___n__q0),
    .stream_s_dout(qw9_vadd_bw__dout),
    .stream_peek_dout(qw9_vadd_bw__dout),
    .stream_s_empty_n(qw9_vadd_bw__empty_n),
    .stream_peek_empty_n(qw9_vadd_bw__empty_n),
    .stream_s_read(qw9_vadd_bw__read),
    .stream_peek_read(),
    .m_axi_mmap_ARADDR(m_axi_rmem9___Stream2Mmap_9___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem9___Stream2Mmap_9___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem9___Stream2Mmap_9___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem9___Stream2Mmap_9___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem9___Stream2Mmap_9___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem9___Stream2Mmap_9___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem9___Stream2Mmap_9___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem9___Stream2Mmap_9___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem9___Stream2Mmap_9___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem9___Stream2Mmap_9___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem9___Stream2Mmap_9___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem9___Stream2Mmap_9___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem9___Stream2Mmap_9___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem9___Stream2Mmap_9___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem9___Stream2Mmap_9___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem9___Stream2Mmap_9___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem9___Stream2Mmap_9___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem9___Stream2Mmap_9___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem9___Stream2Mmap_9___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem9___Stream2Mmap_9___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem9___Stream2Mmap_9___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem9___Stream2Mmap_9___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem9___Stream2Mmap_9___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem9___Stream2Mmap_9___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem9___Stream2Mmap_9___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem9___Stream2Mmap_9___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem9___Stream2Mmap_9___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem9___Stream2Mmap_9___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem9___Stream2Mmap_9___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem9___Stream2Mmap_9___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem9___Stream2Mmap_9___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem9___Stream2Mmap_9___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem9___Stream2Mmap_9___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem9___Stream2Mmap_9___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem9___Stream2Mmap_9___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem9___Stream2Mmap_9___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem9___Stream2Mmap_9___mmap_AWQOS),
    .mmap_offset(Stream2Mmap_9___rmem9__q0)
  );


  (* keep_hierarchy = "yes" *) Stream2Mmap
  Stream2Mmap_10
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Stream2Mmap_10__ap_start),
    .ap_done(Stream2Mmap_10__ap_done),
    .ap_idle(Stream2Mmap_10__ap_idle),
    .ap_ready(Stream2Mmap_10__ap_ready),
    .n(Stream2Mmap_10___n__q0),
    .stream_s_dout(qw10_vadd_bw__dout),
    .stream_peek_dout(qw10_vadd_bw__dout),
    .stream_s_empty_n(qw10_vadd_bw__empty_n),
    .stream_peek_empty_n(qw10_vadd_bw__empty_n),
    .stream_s_read(qw10_vadd_bw__read),
    .stream_peek_read(),
    .m_axi_mmap_ARADDR(m_axi_rmem10___Stream2Mmap_10___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem10___Stream2Mmap_10___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem10___Stream2Mmap_10___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem10___Stream2Mmap_10___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem10___Stream2Mmap_10___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem10___Stream2Mmap_10___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem10___Stream2Mmap_10___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem10___Stream2Mmap_10___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem10___Stream2Mmap_10___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem10___Stream2Mmap_10___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem10___Stream2Mmap_10___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem10___Stream2Mmap_10___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem10___Stream2Mmap_10___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem10___Stream2Mmap_10___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem10___Stream2Mmap_10___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem10___Stream2Mmap_10___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem10___Stream2Mmap_10___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem10___Stream2Mmap_10___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem10___Stream2Mmap_10___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem10___Stream2Mmap_10___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem10___Stream2Mmap_10___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem10___Stream2Mmap_10___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem10___Stream2Mmap_10___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem10___Stream2Mmap_10___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem10___Stream2Mmap_10___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem10___Stream2Mmap_10___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem10___Stream2Mmap_10___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem10___Stream2Mmap_10___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem10___Stream2Mmap_10___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem10___Stream2Mmap_10___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem10___Stream2Mmap_10___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem10___Stream2Mmap_10___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem10___Stream2Mmap_10___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem10___Stream2Mmap_10___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem10___Stream2Mmap_10___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem10___Stream2Mmap_10___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem10___Stream2Mmap_10___mmap_AWQOS),
    .mmap_offset(Stream2Mmap_10___rmem10__q0)
  );


  (* keep_hierarchy = "yes" *) Stream2Mmap
  Stream2Mmap_11
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Stream2Mmap_11__ap_start),
    .ap_done(Stream2Mmap_11__ap_done),
    .ap_idle(Stream2Mmap_11__ap_idle),
    .ap_ready(Stream2Mmap_11__ap_ready),
    .n(Stream2Mmap_11___n__q0),
    .stream_s_dout(qw11_vadd_bw__dout),
    .stream_peek_dout(qw11_vadd_bw__dout),
    .stream_s_empty_n(qw11_vadd_bw__empty_n),
    .stream_peek_empty_n(qw11_vadd_bw__empty_n),
    .stream_s_read(qw11_vadd_bw__read),
    .stream_peek_read(),
    .m_axi_mmap_ARADDR(m_axi_rmem11___Stream2Mmap_11___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem11___Stream2Mmap_11___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem11___Stream2Mmap_11___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem11___Stream2Mmap_11___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem11___Stream2Mmap_11___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem11___Stream2Mmap_11___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem11___Stream2Mmap_11___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem11___Stream2Mmap_11___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem11___Stream2Mmap_11___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem11___Stream2Mmap_11___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem11___Stream2Mmap_11___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem11___Stream2Mmap_11___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem11___Stream2Mmap_11___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem11___Stream2Mmap_11___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem11___Stream2Mmap_11___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem11___Stream2Mmap_11___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem11___Stream2Mmap_11___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem11___Stream2Mmap_11___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem11___Stream2Mmap_11___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem11___Stream2Mmap_11___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem11___Stream2Mmap_11___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem11___Stream2Mmap_11___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem11___Stream2Mmap_11___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem11___Stream2Mmap_11___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem11___Stream2Mmap_11___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem11___Stream2Mmap_11___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem11___Stream2Mmap_11___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem11___Stream2Mmap_11___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem11___Stream2Mmap_11___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem11___Stream2Mmap_11___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem11___Stream2Mmap_11___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem11___Stream2Mmap_11___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem11___Stream2Mmap_11___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem11___Stream2Mmap_11___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem11___Stream2Mmap_11___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem11___Stream2Mmap_11___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem11___Stream2Mmap_11___mmap_AWQOS),
    .mmap_offset(Stream2Mmap_11___rmem11__q0)
  );


  (* keep_hierarchy = "yes" *) Stream2Mmap
  Stream2Mmap_12
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Stream2Mmap_12__ap_start),
    .ap_done(Stream2Mmap_12__ap_done),
    .ap_idle(Stream2Mmap_12__ap_idle),
    .ap_ready(Stream2Mmap_12__ap_ready),
    .n(Stream2Mmap_12___n__q0),
    .stream_s_dout(qw12_vadd_bw__dout),
    .stream_peek_dout(qw12_vadd_bw__dout),
    .stream_s_empty_n(qw12_vadd_bw__empty_n),
    .stream_peek_empty_n(qw12_vadd_bw__empty_n),
    .stream_s_read(qw12_vadd_bw__read),
    .stream_peek_read(),
    .m_axi_mmap_ARADDR(m_axi_rmem12___Stream2Mmap_12___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem12___Stream2Mmap_12___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem12___Stream2Mmap_12___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem12___Stream2Mmap_12___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem12___Stream2Mmap_12___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem12___Stream2Mmap_12___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem12___Stream2Mmap_12___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem12___Stream2Mmap_12___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem12___Stream2Mmap_12___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem12___Stream2Mmap_12___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem12___Stream2Mmap_12___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem12___Stream2Mmap_12___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem12___Stream2Mmap_12___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem12___Stream2Mmap_12___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem12___Stream2Mmap_12___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem12___Stream2Mmap_12___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem12___Stream2Mmap_12___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem12___Stream2Mmap_12___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem12___Stream2Mmap_12___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem12___Stream2Mmap_12___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem12___Stream2Mmap_12___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem12___Stream2Mmap_12___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem12___Stream2Mmap_12___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem12___Stream2Mmap_12___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem12___Stream2Mmap_12___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem12___Stream2Mmap_12___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem12___Stream2Mmap_12___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem12___Stream2Mmap_12___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem12___Stream2Mmap_12___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem12___Stream2Mmap_12___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem12___Stream2Mmap_12___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem12___Stream2Mmap_12___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem12___Stream2Mmap_12___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem12___Stream2Mmap_12___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem12___Stream2Mmap_12___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem12___Stream2Mmap_12___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem12___Stream2Mmap_12___mmap_AWQOS),
    .mmap_offset(Stream2Mmap_12___rmem12__q0)
  );


  (* keep_hierarchy = "yes" *) Stream2Mmap
  Stream2Mmap_13
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Stream2Mmap_13__ap_start),
    .ap_done(Stream2Mmap_13__ap_done),
    .ap_idle(Stream2Mmap_13__ap_idle),
    .ap_ready(Stream2Mmap_13__ap_ready),
    .n(Stream2Mmap_13___n__q0),
    .stream_s_dout(qw13_vadd_bw__dout),
    .stream_peek_dout(qw13_vadd_bw__dout),
    .stream_s_empty_n(qw13_vadd_bw__empty_n),
    .stream_peek_empty_n(qw13_vadd_bw__empty_n),
    .stream_s_read(qw13_vadd_bw__read),
    .stream_peek_read(),
    .m_axi_mmap_ARADDR(m_axi_rmem13___Stream2Mmap_13___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem13___Stream2Mmap_13___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem13___Stream2Mmap_13___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem13___Stream2Mmap_13___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem13___Stream2Mmap_13___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem13___Stream2Mmap_13___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem13___Stream2Mmap_13___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem13___Stream2Mmap_13___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem13___Stream2Mmap_13___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem13___Stream2Mmap_13___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem13___Stream2Mmap_13___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem13___Stream2Mmap_13___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem13___Stream2Mmap_13___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem13___Stream2Mmap_13___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem13___Stream2Mmap_13___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem13___Stream2Mmap_13___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem13___Stream2Mmap_13___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem13___Stream2Mmap_13___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem13___Stream2Mmap_13___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem13___Stream2Mmap_13___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem13___Stream2Mmap_13___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem13___Stream2Mmap_13___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem13___Stream2Mmap_13___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem13___Stream2Mmap_13___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem13___Stream2Mmap_13___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem13___Stream2Mmap_13___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem13___Stream2Mmap_13___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem13___Stream2Mmap_13___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem13___Stream2Mmap_13___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem13___Stream2Mmap_13___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem13___Stream2Mmap_13___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem13___Stream2Mmap_13___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem13___Stream2Mmap_13___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem13___Stream2Mmap_13___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem13___Stream2Mmap_13___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem13___Stream2Mmap_13___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem13___Stream2Mmap_13___mmap_AWQOS),
    .mmap_offset(Stream2Mmap_13___rmem13__q0)
  );


  (* keep_hierarchy = "yes" *) Stream2Mmap
  Stream2Mmap_14
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Stream2Mmap_14__ap_start),
    .ap_done(Stream2Mmap_14__ap_done),
    .ap_idle(Stream2Mmap_14__ap_idle),
    .ap_ready(Stream2Mmap_14__ap_ready),
    .n(Stream2Mmap_14___n__q0),
    .stream_s_dout(qw14_vadd_bw__dout),
    .stream_peek_dout(qw14_vadd_bw__dout),
    .stream_s_empty_n(qw14_vadd_bw__empty_n),
    .stream_peek_empty_n(qw14_vadd_bw__empty_n),
    .stream_s_read(qw14_vadd_bw__read),
    .stream_peek_read(),
    .m_axi_mmap_ARADDR(m_axi_rmem14___Stream2Mmap_14___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem14___Stream2Mmap_14___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem14___Stream2Mmap_14___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem14___Stream2Mmap_14___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem14___Stream2Mmap_14___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem14___Stream2Mmap_14___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem14___Stream2Mmap_14___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem14___Stream2Mmap_14___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem14___Stream2Mmap_14___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem14___Stream2Mmap_14___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem14___Stream2Mmap_14___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem14___Stream2Mmap_14___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem14___Stream2Mmap_14___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem14___Stream2Mmap_14___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem14___Stream2Mmap_14___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem14___Stream2Mmap_14___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem14___Stream2Mmap_14___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem14___Stream2Mmap_14___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem14___Stream2Mmap_14___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem14___Stream2Mmap_14___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem14___Stream2Mmap_14___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem14___Stream2Mmap_14___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem14___Stream2Mmap_14___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem14___Stream2Mmap_14___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem14___Stream2Mmap_14___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem14___Stream2Mmap_14___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem14___Stream2Mmap_14___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem14___Stream2Mmap_14___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem14___Stream2Mmap_14___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem14___Stream2Mmap_14___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem14___Stream2Mmap_14___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem14___Stream2Mmap_14___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem14___Stream2Mmap_14___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem14___Stream2Mmap_14___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem14___Stream2Mmap_14___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem14___Stream2Mmap_14___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem14___Stream2Mmap_14___mmap_AWQOS),
    .mmap_offset(Stream2Mmap_14___rmem14__q0)
  );


  (* keep_hierarchy = "yes" *) Stream2Mmap
  Stream2Mmap_15
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Stream2Mmap_15__ap_start),
    .ap_done(Stream2Mmap_15__ap_done),
    .ap_idle(Stream2Mmap_15__ap_idle),
    .ap_ready(Stream2Mmap_15__ap_ready),
    .n(Stream2Mmap_15___n__q0),
    .stream_s_dout(qw15_vadd_bw__dout),
    .stream_peek_dout(qw15_vadd_bw__dout),
    .stream_s_empty_n(qw15_vadd_bw__empty_n),
    .stream_peek_empty_n(qw15_vadd_bw__empty_n),
    .stream_s_read(qw15_vadd_bw__read),
    .stream_peek_read(),
    .m_axi_mmap_ARADDR(m_axi_rmem15___Stream2Mmap_15___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem15___Stream2Mmap_15___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem15___Stream2Mmap_15___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem15___Stream2Mmap_15___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem15___Stream2Mmap_15___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem15___Stream2Mmap_15___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem15___Stream2Mmap_15___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem15___Stream2Mmap_15___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem15___Stream2Mmap_15___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem15___Stream2Mmap_15___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem15___Stream2Mmap_15___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem15___Stream2Mmap_15___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem15___Stream2Mmap_15___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem15___Stream2Mmap_15___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem15___Stream2Mmap_15___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem15___Stream2Mmap_15___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem15___Stream2Mmap_15___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem15___Stream2Mmap_15___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem15___Stream2Mmap_15___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem15___Stream2Mmap_15___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem15___Stream2Mmap_15___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem15___Stream2Mmap_15___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem15___Stream2Mmap_15___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem15___Stream2Mmap_15___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem15___Stream2Mmap_15___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem15___Stream2Mmap_15___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem15___Stream2Mmap_15___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem15___Stream2Mmap_15___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem15___Stream2Mmap_15___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem15___Stream2Mmap_15___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem15___Stream2Mmap_15___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem15___Stream2Mmap_15___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem15___Stream2Mmap_15___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem15___Stream2Mmap_15___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem15___Stream2Mmap_15___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem15___Stream2Mmap_15___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem15___Stream2Mmap_15___mmap_AWQOS),
    .mmap_offset(Stream2Mmap_15___rmem15__q0)
  );


  (* keep_hierarchy = "yes" *) Stream2Mmap
  Stream2Mmap_16
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Stream2Mmap_16__ap_start),
    .ap_done(Stream2Mmap_16__ap_done),
    .ap_idle(Stream2Mmap_16__ap_idle),
    .ap_ready(Stream2Mmap_16__ap_ready),
    .n(Stream2Mmap_16___n__q0),
    .stream_s_dout(qw16_vadd_bw__dout),
    .stream_peek_dout(qw16_vadd_bw__dout),
    .stream_s_empty_n(qw16_vadd_bw__empty_n),
    .stream_peek_empty_n(qw16_vadd_bw__empty_n),
    .stream_s_read(qw16_vadd_bw__read),
    .stream_peek_read(),
    .m_axi_mmap_ARADDR(m_axi_rmem16___Stream2Mmap_16___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem16___Stream2Mmap_16___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem16___Stream2Mmap_16___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem16___Stream2Mmap_16___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem16___Stream2Mmap_16___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem16___Stream2Mmap_16___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem16___Stream2Mmap_16___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem16___Stream2Mmap_16___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem16___Stream2Mmap_16___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem16___Stream2Mmap_16___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem16___Stream2Mmap_16___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem16___Stream2Mmap_16___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem16___Stream2Mmap_16___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem16___Stream2Mmap_16___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem16___Stream2Mmap_16___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem16___Stream2Mmap_16___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem16___Stream2Mmap_16___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem16___Stream2Mmap_16___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem16___Stream2Mmap_16___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem16___Stream2Mmap_16___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem16___Stream2Mmap_16___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem16___Stream2Mmap_16___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem16___Stream2Mmap_16___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem16___Stream2Mmap_16___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem16___Stream2Mmap_16___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem16___Stream2Mmap_16___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem16___Stream2Mmap_16___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem16___Stream2Mmap_16___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem16___Stream2Mmap_16___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem16___Stream2Mmap_16___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem16___Stream2Mmap_16___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem16___Stream2Mmap_16___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem16___Stream2Mmap_16___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem16___Stream2Mmap_16___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem16___Stream2Mmap_16___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem16___Stream2Mmap_16___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem16___Stream2Mmap_16___mmap_AWQOS),
    .mmap_offset(Stream2Mmap_16___rmem16__q0)
  );


  (* keep_hierarchy = "yes" *) Stream2Mmap
  Stream2Mmap_17
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Stream2Mmap_17__ap_start),
    .ap_done(Stream2Mmap_17__ap_done),
    .ap_idle(Stream2Mmap_17__ap_idle),
    .ap_ready(Stream2Mmap_17__ap_ready),
    .n(Stream2Mmap_17___n__q0),
    .stream_s_dout(qw17_vadd_bw__dout),
    .stream_peek_dout(qw17_vadd_bw__dout),
    .stream_s_empty_n(qw17_vadd_bw__empty_n),
    .stream_peek_empty_n(qw17_vadd_bw__empty_n),
    .stream_s_read(qw17_vadd_bw__read),
    .stream_peek_read(),
    .m_axi_mmap_ARADDR(m_axi_rmem17___Stream2Mmap_17___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem17___Stream2Mmap_17___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem17___Stream2Mmap_17___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem17___Stream2Mmap_17___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem17___Stream2Mmap_17___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem17___Stream2Mmap_17___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem17___Stream2Mmap_17___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem17___Stream2Mmap_17___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem17___Stream2Mmap_17___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem17___Stream2Mmap_17___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem17___Stream2Mmap_17___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem17___Stream2Mmap_17___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem17___Stream2Mmap_17___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem17___Stream2Mmap_17___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem17___Stream2Mmap_17___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem17___Stream2Mmap_17___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem17___Stream2Mmap_17___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem17___Stream2Mmap_17___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem17___Stream2Mmap_17___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem17___Stream2Mmap_17___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem17___Stream2Mmap_17___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem17___Stream2Mmap_17___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem17___Stream2Mmap_17___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem17___Stream2Mmap_17___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem17___Stream2Mmap_17___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem17___Stream2Mmap_17___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem17___Stream2Mmap_17___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem17___Stream2Mmap_17___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem17___Stream2Mmap_17___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem17___Stream2Mmap_17___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem17___Stream2Mmap_17___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem17___Stream2Mmap_17___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem17___Stream2Mmap_17___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem17___Stream2Mmap_17___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem17___Stream2Mmap_17___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem17___Stream2Mmap_17___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem17___Stream2Mmap_17___mmap_AWQOS),
    .mmap_offset(Stream2Mmap_17___rmem17__q0)
  );


  (* keep_hierarchy = "yes" *) Stream2Mmap
  Stream2Mmap_18
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Stream2Mmap_18__ap_start),
    .ap_done(Stream2Mmap_18__ap_done),
    .ap_idle(Stream2Mmap_18__ap_idle),
    .ap_ready(Stream2Mmap_18__ap_ready),
    .n(Stream2Mmap_18___n__q0),
    .stream_s_dout(qw18_vadd_bw__dout),
    .stream_peek_dout(qw18_vadd_bw__dout),
    .stream_s_empty_n(qw18_vadd_bw__empty_n),
    .stream_peek_empty_n(qw18_vadd_bw__empty_n),
    .stream_s_read(qw18_vadd_bw__read),
    .stream_peek_read(),
    .m_axi_mmap_ARADDR(m_axi_rmem18___Stream2Mmap_18___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem18___Stream2Mmap_18___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem18___Stream2Mmap_18___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem18___Stream2Mmap_18___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem18___Stream2Mmap_18___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem18___Stream2Mmap_18___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem18___Stream2Mmap_18___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem18___Stream2Mmap_18___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem18___Stream2Mmap_18___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem18___Stream2Mmap_18___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem18___Stream2Mmap_18___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem18___Stream2Mmap_18___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem18___Stream2Mmap_18___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem18___Stream2Mmap_18___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem18___Stream2Mmap_18___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem18___Stream2Mmap_18___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem18___Stream2Mmap_18___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem18___Stream2Mmap_18___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem18___Stream2Mmap_18___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem18___Stream2Mmap_18___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem18___Stream2Mmap_18___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem18___Stream2Mmap_18___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem18___Stream2Mmap_18___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem18___Stream2Mmap_18___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem18___Stream2Mmap_18___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem18___Stream2Mmap_18___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem18___Stream2Mmap_18___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem18___Stream2Mmap_18___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem18___Stream2Mmap_18___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem18___Stream2Mmap_18___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem18___Stream2Mmap_18___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem18___Stream2Mmap_18___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem18___Stream2Mmap_18___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem18___Stream2Mmap_18___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem18___Stream2Mmap_18___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem18___Stream2Mmap_18___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem18___Stream2Mmap_18___mmap_AWQOS),
    .mmap_offset(Stream2Mmap_18___rmem18__q0)
  );


  (* keep_hierarchy = "yes" *) Stream2Mmap
  Stream2Mmap_19
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Stream2Mmap_19__ap_start),
    .ap_done(Stream2Mmap_19__ap_done),
    .ap_idle(Stream2Mmap_19__ap_idle),
    .ap_ready(Stream2Mmap_19__ap_ready),
    .n(Stream2Mmap_19___n__q0),
    .stream_s_dout(qw19_vadd_bw__dout),
    .stream_peek_dout(qw19_vadd_bw__dout),
    .stream_s_empty_n(qw19_vadd_bw__empty_n),
    .stream_peek_empty_n(qw19_vadd_bw__empty_n),
    .stream_s_read(qw19_vadd_bw__read),
    .stream_peek_read(),
    .m_axi_mmap_ARADDR(m_axi_rmem19___Stream2Mmap_19___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem19___Stream2Mmap_19___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem19___Stream2Mmap_19___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem19___Stream2Mmap_19___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem19___Stream2Mmap_19___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem19___Stream2Mmap_19___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem19___Stream2Mmap_19___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem19___Stream2Mmap_19___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem19___Stream2Mmap_19___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem19___Stream2Mmap_19___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem19___Stream2Mmap_19___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem19___Stream2Mmap_19___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem19___Stream2Mmap_19___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem19___Stream2Mmap_19___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem19___Stream2Mmap_19___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem19___Stream2Mmap_19___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem19___Stream2Mmap_19___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem19___Stream2Mmap_19___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem19___Stream2Mmap_19___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem19___Stream2Mmap_19___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem19___Stream2Mmap_19___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem19___Stream2Mmap_19___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem19___Stream2Mmap_19___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem19___Stream2Mmap_19___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem19___Stream2Mmap_19___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem19___Stream2Mmap_19___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem19___Stream2Mmap_19___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem19___Stream2Mmap_19___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem19___Stream2Mmap_19___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem19___Stream2Mmap_19___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem19___Stream2Mmap_19___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem19___Stream2Mmap_19___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem19___Stream2Mmap_19___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem19___Stream2Mmap_19___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem19___Stream2Mmap_19___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem19___Stream2Mmap_19___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem19___Stream2Mmap_19___mmap_AWQOS),
    .mmap_offset(Stream2Mmap_19___rmem19__q0)
  );


  (* keep_hierarchy = "yes" *) Stream2Mmap
  Stream2Mmap_20
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Stream2Mmap_20__ap_start),
    .ap_done(Stream2Mmap_20__ap_done),
    .ap_idle(Stream2Mmap_20__ap_idle),
    .ap_ready(Stream2Mmap_20__ap_ready),
    .n(Stream2Mmap_20___n__q0),
    .stream_s_dout(qw20_vadd_bw__dout),
    .stream_peek_dout(qw20_vadd_bw__dout),
    .stream_s_empty_n(qw20_vadd_bw__empty_n),
    .stream_peek_empty_n(qw20_vadd_bw__empty_n),
    .stream_s_read(qw20_vadd_bw__read),
    .stream_peek_read(),
    .m_axi_mmap_ARADDR(m_axi_rmem20___Stream2Mmap_20___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem20___Stream2Mmap_20___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem20___Stream2Mmap_20___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem20___Stream2Mmap_20___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem20___Stream2Mmap_20___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem20___Stream2Mmap_20___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem20___Stream2Mmap_20___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem20___Stream2Mmap_20___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem20___Stream2Mmap_20___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem20___Stream2Mmap_20___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem20___Stream2Mmap_20___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem20___Stream2Mmap_20___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem20___Stream2Mmap_20___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem20___Stream2Mmap_20___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem20___Stream2Mmap_20___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem20___Stream2Mmap_20___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem20___Stream2Mmap_20___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem20___Stream2Mmap_20___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem20___Stream2Mmap_20___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem20___Stream2Mmap_20___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem20___Stream2Mmap_20___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem20___Stream2Mmap_20___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem20___Stream2Mmap_20___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem20___Stream2Mmap_20___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem20___Stream2Mmap_20___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem20___Stream2Mmap_20___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem20___Stream2Mmap_20___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem20___Stream2Mmap_20___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem20___Stream2Mmap_20___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem20___Stream2Mmap_20___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem20___Stream2Mmap_20___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem20___Stream2Mmap_20___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem20___Stream2Mmap_20___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem20___Stream2Mmap_20___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem20___Stream2Mmap_20___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem20___Stream2Mmap_20___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem20___Stream2Mmap_20___mmap_AWQOS),
    .mmap_offset(Stream2Mmap_20___rmem20__q0)
  );


  (* keep_hierarchy = "yes" *) Stream2Mmap
  Stream2Mmap_21
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Stream2Mmap_21__ap_start),
    .ap_done(Stream2Mmap_21__ap_done),
    .ap_idle(Stream2Mmap_21__ap_idle),
    .ap_ready(Stream2Mmap_21__ap_ready),
    .n(Stream2Mmap_21___n__q0),
    .stream_s_dout(qw21_vadd_bw__dout),
    .stream_peek_dout(qw21_vadd_bw__dout),
    .stream_s_empty_n(qw21_vadd_bw__empty_n),
    .stream_peek_empty_n(qw21_vadd_bw__empty_n),
    .stream_s_read(qw21_vadd_bw__read),
    .stream_peek_read(),
    .m_axi_mmap_ARADDR(m_axi_rmem21___Stream2Mmap_21___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem21___Stream2Mmap_21___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem21___Stream2Mmap_21___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem21___Stream2Mmap_21___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem21___Stream2Mmap_21___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem21___Stream2Mmap_21___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem21___Stream2Mmap_21___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem21___Stream2Mmap_21___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem21___Stream2Mmap_21___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem21___Stream2Mmap_21___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem21___Stream2Mmap_21___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem21___Stream2Mmap_21___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem21___Stream2Mmap_21___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem21___Stream2Mmap_21___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem21___Stream2Mmap_21___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem21___Stream2Mmap_21___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem21___Stream2Mmap_21___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem21___Stream2Mmap_21___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem21___Stream2Mmap_21___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem21___Stream2Mmap_21___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem21___Stream2Mmap_21___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem21___Stream2Mmap_21___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem21___Stream2Mmap_21___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem21___Stream2Mmap_21___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem21___Stream2Mmap_21___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem21___Stream2Mmap_21___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem21___Stream2Mmap_21___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem21___Stream2Mmap_21___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem21___Stream2Mmap_21___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem21___Stream2Mmap_21___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem21___Stream2Mmap_21___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem21___Stream2Mmap_21___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem21___Stream2Mmap_21___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem21___Stream2Mmap_21___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem21___Stream2Mmap_21___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem21___Stream2Mmap_21___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem21___Stream2Mmap_21___mmap_AWQOS),
    .mmap_offset(Stream2Mmap_21___rmem21__q0)
  );


  (* keep_hierarchy = "yes" *) Stream2Mmap
  Stream2Mmap_22
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Stream2Mmap_22__ap_start),
    .ap_done(Stream2Mmap_22__ap_done),
    .ap_idle(Stream2Mmap_22__ap_idle),
    .ap_ready(Stream2Mmap_22__ap_ready),
    .n(Stream2Mmap_22___n__q0),
    .stream_s_dout(qw22_vadd_bw__dout),
    .stream_peek_dout(qw22_vadd_bw__dout),
    .stream_s_empty_n(qw22_vadd_bw__empty_n),
    .stream_peek_empty_n(qw22_vadd_bw__empty_n),
    .stream_s_read(qw22_vadd_bw__read),
    .stream_peek_read(),
    .m_axi_mmap_ARADDR(m_axi_rmem22___Stream2Mmap_22___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem22___Stream2Mmap_22___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem22___Stream2Mmap_22___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem22___Stream2Mmap_22___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem22___Stream2Mmap_22___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem22___Stream2Mmap_22___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem22___Stream2Mmap_22___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem22___Stream2Mmap_22___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem22___Stream2Mmap_22___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem22___Stream2Mmap_22___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem22___Stream2Mmap_22___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem22___Stream2Mmap_22___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem22___Stream2Mmap_22___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem22___Stream2Mmap_22___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem22___Stream2Mmap_22___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem22___Stream2Mmap_22___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem22___Stream2Mmap_22___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem22___Stream2Mmap_22___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem22___Stream2Mmap_22___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem22___Stream2Mmap_22___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem22___Stream2Mmap_22___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem22___Stream2Mmap_22___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem22___Stream2Mmap_22___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem22___Stream2Mmap_22___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem22___Stream2Mmap_22___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem22___Stream2Mmap_22___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem22___Stream2Mmap_22___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem22___Stream2Mmap_22___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem22___Stream2Mmap_22___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem22___Stream2Mmap_22___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem22___Stream2Mmap_22___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem22___Stream2Mmap_22___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem22___Stream2Mmap_22___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem22___Stream2Mmap_22___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem22___Stream2Mmap_22___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem22___Stream2Mmap_22___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem22___Stream2Mmap_22___mmap_AWQOS),
    .mmap_offset(Stream2Mmap_22___rmem22__q0)
  );


  (* keep_hierarchy = "yes" *) Stream2Mmap
  Stream2Mmap_23
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Stream2Mmap_23__ap_start),
    .ap_done(Stream2Mmap_23__ap_done),
    .ap_idle(Stream2Mmap_23__ap_idle),
    .ap_ready(Stream2Mmap_23__ap_ready),
    .n(Stream2Mmap_23___n__q0),
    .stream_s_dout(qw23_vadd_bw__dout),
    .stream_peek_dout(qw23_vadd_bw__dout),
    .stream_s_empty_n(qw23_vadd_bw__empty_n),
    .stream_peek_empty_n(qw23_vadd_bw__empty_n),
    .stream_s_read(qw23_vadd_bw__read),
    .stream_peek_read(),
    .m_axi_mmap_ARADDR(m_axi_rmem23___Stream2Mmap_23___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem23___Stream2Mmap_23___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem23___Stream2Mmap_23___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem23___Stream2Mmap_23___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem23___Stream2Mmap_23___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem23___Stream2Mmap_23___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem23___Stream2Mmap_23___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem23___Stream2Mmap_23___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem23___Stream2Mmap_23___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem23___Stream2Mmap_23___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem23___Stream2Mmap_23___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem23___Stream2Mmap_23___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem23___Stream2Mmap_23___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem23___Stream2Mmap_23___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem23___Stream2Mmap_23___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem23___Stream2Mmap_23___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem23___Stream2Mmap_23___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem23___Stream2Mmap_23___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem23___Stream2Mmap_23___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem23___Stream2Mmap_23___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem23___Stream2Mmap_23___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem23___Stream2Mmap_23___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem23___Stream2Mmap_23___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem23___Stream2Mmap_23___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem23___Stream2Mmap_23___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem23___Stream2Mmap_23___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem23___Stream2Mmap_23___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem23___Stream2Mmap_23___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem23___Stream2Mmap_23___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem23___Stream2Mmap_23___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem23___Stream2Mmap_23___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem23___Stream2Mmap_23___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem23___Stream2Mmap_23___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem23___Stream2Mmap_23___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem23___Stream2Mmap_23___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem23___Stream2Mmap_23___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem23___Stream2Mmap_23___mmap_AWQOS),
    .mmap_offset(Stream2Mmap_23___rmem23__q0)
  );


  (* keep_hierarchy = "yes" *) Stream2Mmap
  Stream2Mmap_24
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Stream2Mmap_24__ap_start),
    .ap_done(Stream2Mmap_24__ap_done),
    .ap_idle(Stream2Mmap_24__ap_idle),
    .ap_ready(Stream2Mmap_24__ap_ready),
    .n(Stream2Mmap_24___n__q0),
    .stream_s_dout(qw24_vadd_bw__dout),
    .stream_peek_dout(qw24_vadd_bw__dout),
    .stream_s_empty_n(qw24_vadd_bw__empty_n),
    .stream_peek_empty_n(qw24_vadd_bw__empty_n),
    .stream_s_read(qw24_vadd_bw__read),
    .stream_peek_read(),
    .m_axi_mmap_ARADDR(m_axi_rmem24___Stream2Mmap_24___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem24___Stream2Mmap_24___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem24___Stream2Mmap_24___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem24___Stream2Mmap_24___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem24___Stream2Mmap_24___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem24___Stream2Mmap_24___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem24___Stream2Mmap_24___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem24___Stream2Mmap_24___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem24___Stream2Mmap_24___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem24___Stream2Mmap_24___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem24___Stream2Mmap_24___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem24___Stream2Mmap_24___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem24___Stream2Mmap_24___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem24___Stream2Mmap_24___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem24___Stream2Mmap_24___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem24___Stream2Mmap_24___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem24___Stream2Mmap_24___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem24___Stream2Mmap_24___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem24___Stream2Mmap_24___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem24___Stream2Mmap_24___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem24___Stream2Mmap_24___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem24___Stream2Mmap_24___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem24___Stream2Mmap_24___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem24___Stream2Mmap_24___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem24___Stream2Mmap_24___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem24___Stream2Mmap_24___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem24___Stream2Mmap_24___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem24___Stream2Mmap_24___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem24___Stream2Mmap_24___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem24___Stream2Mmap_24___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem24___Stream2Mmap_24___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem24___Stream2Mmap_24___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem24___Stream2Mmap_24___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem24___Stream2Mmap_24___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem24___Stream2Mmap_24___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem24___Stream2Mmap_24___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem24___Stream2Mmap_24___mmap_AWQOS),
    .mmap_offset(Stream2Mmap_24___rmem24__q0)
  );


  (* keep_hierarchy = "yes" *) Stream2Mmap
  Stream2Mmap_25
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Stream2Mmap_25__ap_start),
    .ap_done(Stream2Mmap_25__ap_done),
    .ap_idle(Stream2Mmap_25__ap_idle),
    .ap_ready(Stream2Mmap_25__ap_ready),
    .n(Stream2Mmap_25___n__q0),
    .stream_s_dout(qw25_vadd_bw__dout),
    .stream_peek_dout(qw25_vadd_bw__dout),
    .stream_s_empty_n(qw25_vadd_bw__empty_n),
    .stream_peek_empty_n(qw25_vadd_bw__empty_n),
    .stream_s_read(qw25_vadd_bw__read),
    .stream_peek_read(),
    .m_axi_mmap_ARADDR(m_axi_rmem25___Stream2Mmap_25___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem25___Stream2Mmap_25___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem25___Stream2Mmap_25___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem25___Stream2Mmap_25___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem25___Stream2Mmap_25___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem25___Stream2Mmap_25___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem25___Stream2Mmap_25___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem25___Stream2Mmap_25___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem25___Stream2Mmap_25___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem25___Stream2Mmap_25___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem25___Stream2Mmap_25___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem25___Stream2Mmap_25___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem25___Stream2Mmap_25___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem25___Stream2Mmap_25___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem25___Stream2Mmap_25___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem25___Stream2Mmap_25___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem25___Stream2Mmap_25___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem25___Stream2Mmap_25___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem25___Stream2Mmap_25___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem25___Stream2Mmap_25___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem25___Stream2Mmap_25___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem25___Stream2Mmap_25___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem25___Stream2Mmap_25___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem25___Stream2Mmap_25___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem25___Stream2Mmap_25___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem25___Stream2Mmap_25___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem25___Stream2Mmap_25___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem25___Stream2Mmap_25___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem25___Stream2Mmap_25___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem25___Stream2Mmap_25___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem25___Stream2Mmap_25___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem25___Stream2Mmap_25___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem25___Stream2Mmap_25___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem25___Stream2Mmap_25___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem25___Stream2Mmap_25___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem25___Stream2Mmap_25___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem25___Stream2Mmap_25___mmap_AWQOS),
    .mmap_offset(Stream2Mmap_25___rmem25__q0)
  );


  (* keep_hierarchy = "yes" *) Stream2Mmap
  Stream2Mmap_26
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Stream2Mmap_26__ap_start),
    .ap_done(Stream2Mmap_26__ap_done),
    .ap_idle(Stream2Mmap_26__ap_idle),
    .ap_ready(Stream2Mmap_26__ap_ready),
    .n(Stream2Mmap_26___n__q0),
    .stream_s_dout(qw26_vadd_bw__dout),
    .stream_peek_dout(qw26_vadd_bw__dout),
    .stream_s_empty_n(qw26_vadd_bw__empty_n),
    .stream_peek_empty_n(qw26_vadd_bw__empty_n),
    .stream_s_read(qw26_vadd_bw__read),
    .stream_peek_read(),
    .m_axi_mmap_ARADDR(m_axi_rmem26___Stream2Mmap_26___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem26___Stream2Mmap_26___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem26___Stream2Mmap_26___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem26___Stream2Mmap_26___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem26___Stream2Mmap_26___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem26___Stream2Mmap_26___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem26___Stream2Mmap_26___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem26___Stream2Mmap_26___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem26___Stream2Mmap_26___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem26___Stream2Mmap_26___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem26___Stream2Mmap_26___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem26___Stream2Mmap_26___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem26___Stream2Mmap_26___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem26___Stream2Mmap_26___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem26___Stream2Mmap_26___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem26___Stream2Mmap_26___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem26___Stream2Mmap_26___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem26___Stream2Mmap_26___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem26___Stream2Mmap_26___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem26___Stream2Mmap_26___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem26___Stream2Mmap_26___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem26___Stream2Mmap_26___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem26___Stream2Mmap_26___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem26___Stream2Mmap_26___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem26___Stream2Mmap_26___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem26___Stream2Mmap_26___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem26___Stream2Mmap_26___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem26___Stream2Mmap_26___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem26___Stream2Mmap_26___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem26___Stream2Mmap_26___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem26___Stream2Mmap_26___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem26___Stream2Mmap_26___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem26___Stream2Mmap_26___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem26___Stream2Mmap_26___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem26___Stream2Mmap_26___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem26___Stream2Mmap_26___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem26___Stream2Mmap_26___mmap_AWQOS),
    .mmap_offset(Stream2Mmap_26___rmem26__q0)
  );


  (* keep_hierarchy = "yes" *) Stream2Mmap
  Stream2Mmap_27
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Stream2Mmap_27__ap_start),
    .ap_done(Stream2Mmap_27__ap_done),
    .ap_idle(Stream2Mmap_27__ap_idle),
    .ap_ready(Stream2Mmap_27__ap_ready),
    .n(Stream2Mmap_27___n__q0),
    .stream_s_dout(qw27_vadd_bw__dout),
    .stream_peek_dout(qw27_vadd_bw__dout),
    .stream_s_empty_n(qw27_vadd_bw__empty_n),
    .stream_peek_empty_n(qw27_vadd_bw__empty_n),
    .stream_s_read(qw27_vadd_bw__read),
    .stream_peek_read(),
    .m_axi_mmap_ARADDR(m_axi_rmem27___Stream2Mmap_27___mmap_ARADDR),
    .m_axi_mmap_ARBURST(m_axi_rmem27___Stream2Mmap_27___mmap_ARBURST),
    .m_axi_mmap_ARID(m_axi_rmem27___Stream2Mmap_27___mmap_ARID),
    .m_axi_mmap_ARLEN(m_axi_rmem27___Stream2Mmap_27___mmap_ARLEN),
    .m_axi_mmap_ARREADY(m_axi_rmem27___Stream2Mmap_27___mmap_ARREADY),
    .m_axi_mmap_ARSIZE(m_axi_rmem27___Stream2Mmap_27___mmap_ARSIZE),
    .m_axi_mmap_ARVALID(m_axi_rmem27___Stream2Mmap_27___mmap_ARVALID),
    .m_axi_mmap_AWADDR(m_axi_rmem27___Stream2Mmap_27___mmap_AWADDR),
    .m_axi_mmap_AWBURST(m_axi_rmem27___Stream2Mmap_27___mmap_AWBURST),
    .m_axi_mmap_AWID(m_axi_rmem27___Stream2Mmap_27___mmap_AWID),
    .m_axi_mmap_AWLEN(m_axi_rmem27___Stream2Mmap_27___mmap_AWLEN),
    .m_axi_mmap_AWREADY(m_axi_rmem27___Stream2Mmap_27___mmap_AWREADY),
    .m_axi_mmap_AWSIZE(m_axi_rmem27___Stream2Mmap_27___mmap_AWSIZE),
    .m_axi_mmap_AWVALID(m_axi_rmem27___Stream2Mmap_27___mmap_AWVALID),
    .m_axi_mmap_BID(m_axi_rmem27___Stream2Mmap_27___mmap_BID),
    .m_axi_mmap_BREADY(m_axi_rmem27___Stream2Mmap_27___mmap_BREADY),
    .m_axi_mmap_BRESP(m_axi_rmem27___Stream2Mmap_27___mmap_BRESP),
    .m_axi_mmap_BVALID(m_axi_rmem27___Stream2Mmap_27___mmap_BVALID),
    .m_axi_mmap_RDATA(m_axi_rmem27___Stream2Mmap_27___mmap_RDATA),
    .m_axi_mmap_RID(m_axi_rmem27___Stream2Mmap_27___mmap_RID),
    .m_axi_mmap_RLAST(m_axi_rmem27___Stream2Mmap_27___mmap_RLAST),
    .m_axi_mmap_RREADY(m_axi_rmem27___Stream2Mmap_27___mmap_RREADY),
    .m_axi_mmap_RRESP(m_axi_rmem27___Stream2Mmap_27___mmap_RRESP),
    .m_axi_mmap_RVALID(m_axi_rmem27___Stream2Mmap_27___mmap_RVALID),
    .m_axi_mmap_WDATA(m_axi_rmem27___Stream2Mmap_27___mmap_WDATA),
    .m_axi_mmap_WLAST(m_axi_rmem27___Stream2Mmap_27___mmap_WLAST),
    .m_axi_mmap_WREADY(m_axi_rmem27___Stream2Mmap_27___mmap_WREADY),
    .m_axi_mmap_WSTRB(m_axi_rmem27___Stream2Mmap_27___mmap_WSTRB),
    .m_axi_mmap_WVALID(m_axi_rmem27___Stream2Mmap_27___mmap_WVALID),
    .m_axi_mmap_ARLOCK(m_axi_rmem27___Stream2Mmap_27___mmap_ARLOCK),
    .m_axi_mmap_ARPROT(m_axi_rmem27___Stream2Mmap_27___mmap_ARPROT),
    .m_axi_mmap_ARQOS(m_axi_rmem27___Stream2Mmap_27___mmap_ARQOS),
    .m_axi_mmap_ARCACHE(m_axi_rmem27___Stream2Mmap_27___mmap_ARCACHE),
    .m_axi_mmap_AWCACHE(m_axi_rmem27___Stream2Mmap_27___mmap_AWCACHE),
    .m_axi_mmap_AWLOCK(m_axi_rmem27___Stream2Mmap_27___mmap_AWLOCK),
    .m_axi_mmap_AWPROT(m_axi_rmem27___Stream2Mmap_27___mmap_AWPROT),
    .m_axi_mmap_AWQOS(m_axi_rmem27___Stream2Mmap_27___mmap_AWQOS),
    .mmap_offset(Stream2Mmap_27___rmem27__q0)
  );


  (* keep_hierarchy = "yes" *) yshift
  yshift_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(yshift_0__ap_start),
    .ap_done(yshift_0__ap_done),
    .ap_idle(yshift_0__ap_idle),
    .ap_ready(yshift_0__ap_ready),
    .n(yshift_0___n__q0),
    .a_s_dout(qr0_vadd_bw__dout),
    .a_peek_dout(qr0_vadd_bw__dout),
    .a_s_empty_n(qr0_vadd_bw__empty_n),
    .a_peek_empty_n(qr0_vadd_bw__empty_n),
    .a_s_read(qr0_vadd_bw__read),
    .a_peek_read(),
    .b_din(qw0_vadd_bw__din),
    .b_full_n(qw0_vadd_bw__full_n),
    .b_write(qw0_vadd_bw__write)
  );


  (* keep_hierarchy = "yes" *) yshift
  yshift_1
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(yshift_1__ap_start),
    .ap_done(yshift_1__ap_done),
    .ap_idle(yshift_1__ap_idle),
    .ap_ready(yshift_1__ap_ready),
    .n(yshift_1___n__q0),
    .a_s_dout(qr1_vadd_bw__dout),
    .a_peek_dout(qr1_vadd_bw__dout),
    .a_s_empty_n(qr1_vadd_bw__empty_n),
    .a_peek_empty_n(qr1_vadd_bw__empty_n),
    .a_s_read(qr1_vadd_bw__read),
    .a_peek_read(),
    .b_din(qw1_vadd_bw__din),
    .b_full_n(qw1_vadd_bw__full_n),
    .b_write(qw1_vadd_bw__write)
  );


  (* keep_hierarchy = "yes" *) yshift
  yshift_2
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(yshift_2__ap_start),
    .ap_done(yshift_2__ap_done),
    .ap_idle(yshift_2__ap_idle),
    .ap_ready(yshift_2__ap_ready),
    .n(yshift_2___n__q0),
    .a_s_dout(qr2_vadd_bw__dout),
    .a_peek_dout(qr2_vadd_bw__dout),
    .a_s_empty_n(qr2_vadd_bw__empty_n),
    .a_peek_empty_n(qr2_vadd_bw__empty_n),
    .a_s_read(qr2_vadd_bw__read),
    .a_peek_read(),
    .b_din(qw2_vadd_bw__din),
    .b_full_n(qw2_vadd_bw__full_n),
    .b_write(qw2_vadd_bw__write)
  );


  (* keep_hierarchy = "yes" *) yshift
  yshift_3
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(yshift_3__ap_start),
    .ap_done(yshift_3__ap_done),
    .ap_idle(yshift_3__ap_idle),
    .ap_ready(yshift_3__ap_ready),
    .n(yshift_3___n__q0),
    .a_s_dout(qr3_vadd_bw__dout),
    .a_peek_dout(qr3_vadd_bw__dout),
    .a_s_empty_n(qr3_vadd_bw__empty_n),
    .a_peek_empty_n(qr3_vadd_bw__empty_n),
    .a_s_read(qr3_vadd_bw__read),
    .a_peek_read(),
    .b_din(qw3_vadd_bw__din),
    .b_full_n(qw3_vadd_bw__full_n),
    .b_write(qw3_vadd_bw__write)
  );


  (* keep_hierarchy = "yes" *) yshift
  yshift_4
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(yshift_4__ap_start),
    .ap_done(yshift_4__ap_done),
    .ap_idle(yshift_4__ap_idle),
    .ap_ready(yshift_4__ap_ready),
    .n(yshift_4___n__q0),
    .a_s_dout(qr4_vadd_bw__dout),
    .a_peek_dout(qr4_vadd_bw__dout),
    .a_s_empty_n(qr4_vadd_bw__empty_n),
    .a_peek_empty_n(qr4_vadd_bw__empty_n),
    .a_s_read(qr4_vadd_bw__read),
    .a_peek_read(),
    .b_din(qw4_vadd_bw__din),
    .b_full_n(qw4_vadd_bw__full_n),
    .b_write(qw4_vadd_bw__write)
  );


  (* keep_hierarchy = "yes" *) yshift
  yshift_5
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(yshift_5__ap_start),
    .ap_done(yshift_5__ap_done),
    .ap_idle(yshift_5__ap_idle),
    .ap_ready(yshift_5__ap_ready),
    .n(yshift_5___n__q0),
    .a_s_dout(qr5_vadd_bw__dout),
    .a_peek_dout(qr5_vadd_bw__dout),
    .a_s_empty_n(qr5_vadd_bw__empty_n),
    .a_peek_empty_n(qr5_vadd_bw__empty_n),
    .a_s_read(qr5_vadd_bw__read),
    .a_peek_read(),
    .b_din(qw5_vadd_bw__din),
    .b_full_n(qw5_vadd_bw__full_n),
    .b_write(qw5_vadd_bw__write)
  );


  (* keep_hierarchy = "yes" *) yshift
  yshift_6
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(yshift_6__ap_start),
    .ap_done(yshift_6__ap_done),
    .ap_idle(yshift_6__ap_idle),
    .ap_ready(yshift_6__ap_ready),
    .n(yshift_6___n__q0),
    .a_s_dout(qr6_vadd_bw__dout),
    .a_peek_dout(qr6_vadd_bw__dout),
    .a_s_empty_n(qr6_vadd_bw__empty_n),
    .a_peek_empty_n(qr6_vadd_bw__empty_n),
    .a_s_read(qr6_vadd_bw__read),
    .a_peek_read(),
    .b_din(qw6_vadd_bw__din),
    .b_full_n(qw6_vadd_bw__full_n),
    .b_write(qw6_vadd_bw__write)
  );


  (* keep_hierarchy = "yes" *) yshift
  yshift_7
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(yshift_7__ap_start),
    .ap_done(yshift_7__ap_done),
    .ap_idle(yshift_7__ap_idle),
    .ap_ready(yshift_7__ap_ready),
    .n(yshift_7___n__q0),
    .a_s_dout(qr7_vadd_bw__dout),
    .a_peek_dout(qr7_vadd_bw__dout),
    .a_s_empty_n(qr7_vadd_bw__empty_n),
    .a_peek_empty_n(qr7_vadd_bw__empty_n),
    .a_s_read(qr7_vadd_bw__read),
    .a_peek_read(),
    .b_din(qw7_vadd_bw__din),
    .b_full_n(qw7_vadd_bw__full_n),
    .b_write(qw7_vadd_bw__write)
  );


  (* keep_hierarchy = "yes" *) yshift
  yshift_8
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(yshift_8__ap_start),
    .ap_done(yshift_8__ap_done),
    .ap_idle(yshift_8__ap_idle),
    .ap_ready(yshift_8__ap_ready),
    .n(yshift_8___n__q0),
    .a_s_dout(qr8_vadd_bw__dout),
    .a_peek_dout(qr8_vadd_bw__dout),
    .a_s_empty_n(qr8_vadd_bw__empty_n),
    .a_peek_empty_n(qr8_vadd_bw__empty_n),
    .a_s_read(qr8_vadd_bw__read),
    .a_peek_read(),
    .b_din(qw8_vadd_bw__din),
    .b_full_n(qw8_vadd_bw__full_n),
    .b_write(qw8_vadd_bw__write)
  );


  (* keep_hierarchy = "yes" *) yshift
  yshift_9
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(yshift_9__ap_start),
    .ap_done(yshift_9__ap_done),
    .ap_idle(yshift_9__ap_idle),
    .ap_ready(yshift_9__ap_ready),
    .n(yshift_9___n__q0),
    .a_s_dout(qr9_vadd_bw__dout),
    .a_peek_dout(qr9_vadd_bw__dout),
    .a_s_empty_n(qr9_vadd_bw__empty_n),
    .a_peek_empty_n(qr9_vadd_bw__empty_n),
    .a_s_read(qr9_vadd_bw__read),
    .a_peek_read(),
    .b_din(qw9_vadd_bw__din),
    .b_full_n(qw9_vadd_bw__full_n),
    .b_write(qw9_vadd_bw__write)
  );


  (* keep_hierarchy = "yes" *) yshift
  yshift_10
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(yshift_10__ap_start),
    .ap_done(yshift_10__ap_done),
    .ap_idle(yshift_10__ap_idle),
    .ap_ready(yshift_10__ap_ready),
    .n(yshift_10___n__q0),
    .a_s_dout(qr10_vadd_bw__dout),
    .a_peek_dout(qr10_vadd_bw__dout),
    .a_s_empty_n(qr10_vadd_bw__empty_n),
    .a_peek_empty_n(qr10_vadd_bw__empty_n),
    .a_s_read(qr10_vadd_bw__read),
    .a_peek_read(),
    .b_din(qw10_vadd_bw__din),
    .b_full_n(qw10_vadd_bw__full_n),
    .b_write(qw10_vadd_bw__write)
  );


  (* keep_hierarchy = "yes" *) yshift
  yshift_11
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(yshift_11__ap_start),
    .ap_done(yshift_11__ap_done),
    .ap_idle(yshift_11__ap_idle),
    .ap_ready(yshift_11__ap_ready),
    .n(yshift_11___n__q0),
    .a_s_dout(qr11_vadd_bw__dout),
    .a_peek_dout(qr11_vadd_bw__dout),
    .a_s_empty_n(qr11_vadd_bw__empty_n),
    .a_peek_empty_n(qr11_vadd_bw__empty_n),
    .a_s_read(qr11_vadd_bw__read),
    .a_peek_read(),
    .b_din(qw11_vadd_bw__din),
    .b_full_n(qw11_vadd_bw__full_n),
    .b_write(qw11_vadd_bw__write)
  );


  (* keep_hierarchy = "yes" *) yshift
  yshift_12
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(yshift_12__ap_start),
    .ap_done(yshift_12__ap_done),
    .ap_idle(yshift_12__ap_idle),
    .ap_ready(yshift_12__ap_ready),
    .n(yshift_12___n__q0),
    .a_s_dout(qr12_vadd_bw__dout),
    .a_peek_dout(qr12_vadd_bw__dout),
    .a_s_empty_n(qr12_vadd_bw__empty_n),
    .a_peek_empty_n(qr12_vadd_bw__empty_n),
    .a_s_read(qr12_vadd_bw__read),
    .a_peek_read(),
    .b_din(qw12_vadd_bw__din),
    .b_full_n(qw12_vadd_bw__full_n),
    .b_write(qw12_vadd_bw__write)
  );


  (* keep_hierarchy = "yes" *) yshift
  yshift_13
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(yshift_13__ap_start),
    .ap_done(yshift_13__ap_done),
    .ap_idle(yshift_13__ap_idle),
    .ap_ready(yshift_13__ap_ready),
    .n(yshift_13___n__q0),
    .a_s_dout(qr13_vadd_bw__dout),
    .a_peek_dout(qr13_vadd_bw__dout),
    .a_s_empty_n(qr13_vadd_bw__empty_n),
    .a_peek_empty_n(qr13_vadd_bw__empty_n),
    .a_s_read(qr13_vadd_bw__read),
    .a_peek_read(),
    .b_din(qw13_vadd_bw__din),
    .b_full_n(qw13_vadd_bw__full_n),
    .b_write(qw13_vadd_bw__write)
  );


  (* keep_hierarchy = "yes" *) yshift
  yshift_14
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(yshift_14__ap_start),
    .ap_done(yshift_14__ap_done),
    .ap_idle(yshift_14__ap_idle),
    .ap_ready(yshift_14__ap_ready),
    .n(yshift_14___n__q0),
    .a_s_dout(qr14_vadd_bw__dout),
    .a_peek_dout(qr14_vadd_bw__dout),
    .a_s_empty_n(qr14_vadd_bw__empty_n),
    .a_peek_empty_n(qr14_vadd_bw__empty_n),
    .a_s_read(qr14_vadd_bw__read),
    .a_peek_read(),
    .b_din(qw14_vadd_bw__din),
    .b_full_n(qw14_vadd_bw__full_n),
    .b_write(qw14_vadd_bw__write)
  );


  (* keep_hierarchy = "yes" *) yshift
  yshift_15
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(yshift_15__ap_start),
    .ap_done(yshift_15__ap_done),
    .ap_idle(yshift_15__ap_idle),
    .ap_ready(yshift_15__ap_ready),
    .n(yshift_15___n__q0),
    .a_s_dout(qr15_vadd_bw__dout),
    .a_peek_dout(qr15_vadd_bw__dout),
    .a_s_empty_n(qr15_vadd_bw__empty_n),
    .a_peek_empty_n(qr15_vadd_bw__empty_n),
    .a_s_read(qr15_vadd_bw__read),
    .a_peek_read(),
    .b_din(qw15_vadd_bw__din),
    .b_full_n(qw15_vadd_bw__full_n),
    .b_write(qw15_vadd_bw__write)
  );


  (* keep_hierarchy = "yes" *) yshift
  yshift_16
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(yshift_16__ap_start),
    .ap_done(yshift_16__ap_done),
    .ap_idle(yshift_16__ap_idle),
    .ap_ready(yshift_16__ap_ready),
    .n(yshift_16___n__q0),
    .a_s_dout(qr16_vadd_bw__dout),
    .a_peek_dout(qr16_vadd_bw__dout),
    .a_s_empty_n(qr16_vadd_bw__empty_n),
    .a_peek_empty_n(qr16_vadd_bw__empty_n),
    .a_s_read(qr16_vadd_bw__read),
    .a_peek_read(),
    .b_din(qw16_vadd_bw__din),
    .b_full_n(qw16_vadd_bw__full_n),
    .b_write(qw16_vadd_bw__write)
  );


  (* keep_hierarchy = "yes" *) yshift
  yshift_17
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(yshift_17__ap_start),
    .ap_done(yshift_17__ap_done),
    .ap_idle(yshift_17__ap_idle),
    .ap_ready(yshift_17__ap_ready),
    .n(yshift_17___n__q0),
    .a_s_dout(qr17_vadd_bw__dout),
    .a_peek_dout(qr17_vadd_bw__dout),
    .a_s_empty_n(qr17_vadd_bw__empty_n),
    .a_peek_empty_n(qr17_vadd_bw__empty_n),
    .a_s_read(qr17_vadd_bw__read),
    .a_peek_read(),
    .b_din(qw17_vadd_bw__din),
    .b_full_n(qw17_vadd_bw__full_n),
    .b_write(qw17_vadd_bw__write)
  );


  (* keep_hierarchy = "yes" *) yshift
  yshift_18
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(yshift_18__ap_start),
    .ap_done(yshift_18__ap_done),
    .ap_idle(yshift_18__ap_idle),
    .ap_ready(yshift_18__ap_ready),
    .n(yshift_18___n__q0),
    .a_s_dout(qr18_vadd_bw__dout),
    .a_peek_dout(qr18_vadd_bw__dout),
    .a_s_empty_n(qr18_vadd_bw__empty_n),
    .a_peek_empty_n(qr18_vadd_bw__empty_n),
    .a_s_read(qr18_vadd_bw__read),
    .a_peek_read(),
    .b_din(qw18_vadd_bw__din),
    .b_full_n(qw18_vadd_bw__full_n),
    .b_write(qw18_vadd_bw__write)
  );


  (* keep_hierarchy = "yes" *) yshift
  yshift_19
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(yshift_19__ap_start),
    .ap_done(yshift_19__ap_done),
    .ap_idle(yshift_19__ap_idle),
    .ap_ready(yshift_19__ap_ready),
    .n(yshift_19___n__q0),
    .a_s_dout(qr19_vadd_bw__dout),
    .a_peek_dout(qr19_vadd_bw__dout),
    .a_s_empty_n(qr19_vadd_bw__empty_n),
    .a_peek_empty_n(qr19_vadd_bw__empty_n),
    .a_s_read(qr19_vadd_bw__read),
    .a_peek_read(),
    .b_din(qw19_vadd_bw__din),
    .b_full_n(qw19_vadd_bw__full_n),
    .b_write(qw19_vadd_bw__write)
  );


  (* keep_hierarchy = "yes" *) yshift
  yshift_20
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(yshift_20__ap_start),
    .ap_done(yshift_20__ap_done),
    .ap_idle(yshift_20__ap_idle),
    .ap_ready(yshift_20__ap_ready),
    .n(yshift_20___n__q0),
    .a_s_dout(qr20_vadd_bw__dout),
    .a_peek_dout(qr20_vadd_bw__dout),
    .a_s_empty_n(qr20_vadd_bw__empty_n),
    .a_peek_empty_n(qr20_vadd_bw__empty_n),
    .a_s_read(qr20_vadd_bw__read),
    .a_peek_read(),
    .b_din(qw20_vadd_bw__din),
    .b_full_n(qw20_vadd_bw__full_n),
    .b_write(qw20_vadd_bw__write)
  );


  (* keep_hierarchy = "yes" *) yshift
  yshift_21
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(yshift_21__ap_start),
    .ap_done(yshift_21__ap_done),
    .ap_idle(yshift_21__ap_idle),
    .ap_ready(yshift_21__ap_ready),
    .n(yshift_21___n__q0),
    .a_s_dout(qr21_vadd_bw__dout),
    .a_peek_dout(qr21_vadd_bw__dout),
    .a_s_empty_n(qr21_vadd_bw__empty_n),
    .a_peek_empty_n(qr21_vadd_bw__empty_n),
    .a_s_read(qr21_vadd_bw__read),
    .a_peek_read(),
    .b_din(qw21_vadd_bw__din),
    .b_full_n(qw21_vadd_bw__full_n),
    .b_write(qw21_vadd_bw__write)
  );


  (* keep_hierarchy = "yes" *) yshift
  yshift_22
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(yshift_22__ap_start),
    .ap_done(yshift_22__ap_done),
    .ap_idle(yshift_22__ap_idle),
    .ap_ready(yshift_22__ap_ready),
    .n(yshift_22___n__q0),
    .a_s_dout(qr22_vadd_bw__dout),
    .a_peek_dout(qr22_vadd_bw__dout),
    .a_s_empty_n(qr22_vadd_bw__empty_n),
    .a_peek_empty_n(qr22_vadd_bw__empty_n),
    .a_s_read(qr22_vadd_bw__read),
    .a_peek_read(),
    .b_din(qw22_vadd_bw__din),
    .b_full_n(qw22_vadd_bw__full_n),
    .b_write(qw22_vadd_bw__write)
  );


  (* keep_hierarchy = "yes" *) yshift
  yshift_23
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(yshift_23__ap_start),
    .ap_done(yshift_23__ap_done),
    .ap_idle(yshift_23__ap_idle),
    .ap_ready(yshift_23__ap_ready),
    .n(yshift_23___n__q0),
    .a_s_dout(qr23_vadd_bw__dout),
    .a_peek_dout(qr23_vadd_bw__dout),
    .a_s_empty_n(qr23_vadd_bw__empty_n),
    .a_peek_empty_n(qr23_vadd_bw__empty_n),
    .a_s_read(qr23_vadd_bw__read),
    .a_peek_read(),
    .b_din(qw23_vadd_bw__din),
    .b_full_n(qw23_vadd_bw__full_n),
    .b_write(qw23_vadd_bw__write)
  );


  (* keep_hierarchy = "yes" *) yshift
  yshift_24
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(yshift_24__ap_start),
    .ap_done(yshift_24__ap_done),
    .ap_idle(yshift_24__ap_idle),
    .ap_ready(yshift_24__ap_ready),
    .n(yshift_24___n__q0),
    .a_s_dout(qr24_vadd_bw__dout),
    .a_peek_dout(qr24_vadd_bw__dout),
    .a_s_empty_n(qr24_vadd_bw__empty_n),
    .a_peek_empty_n(qr24_vadd_bw__empty_n),
    .a_s_read(qr24_vadd_bw__read),
    .a_peek_read(),
    .b_din(qw24_vadd_bw__din),
    .b_full_n(qw24_vadd_bw__full_n),
    .b_write(qw24_vadd_bw__write)
  );


  (* keep_hierarchy = "yes" *) yshift
  yshift_25
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(yshift_25__ap_start),
    .ap_done(yshift_25__ap_done),
    .ap_idle(yshift_25__ap_idle),
    .ap_ready(yshift_25__ap_ready),
    .n(yshift_25___n__q0),
    .a_s_dout(qr25_vadd_bw__dout),
    .a_peek_dout(qr25_vadd_bw__dout),
    .a_s_empty_n(qr25_vadd_bw__empty_n),
    .a_peek_empty_n(qr25_vadd_bw__empty_n),
    .a_s_read(qr25_vadd_bw__read),
    .a_peek_read(),
    .b_din(qw25_vadd_bw__din),
    .b_full_n(qw25_vadd_bw__full_n),
    .b_write(qw25_vadd_bw__write)
  );


  (* keep_hierarchy = "yes" *) yshift
  yshift_26
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(yshift_26__ap_start),
    .ap_done(yshift_26__ap_done),
    .ap_idle(yshift_26__ap_idle),
    .ap_ready(yshift_26__ap_ready),
    .n(yshift_26___n__q0),
    .a_s_dout(qr26_vadd_bw__dout),
    .a_peek_dout(qr26_vadd_bw__dout),
    .a_s_empty_n(qr26_vadd_bw__empty_n),
    .a_peek_empty_n(qr26_vadd_bw__empty_n),
    .a_s_read(qr26_vadd_bw__read),
    .a_peek_read(),
    .b_din(qw26_vadd_bw__din),
    .b_full_n(qw26_vadd_bw__full_n),
    .b_write(qw26_vadd_bw__write)
  );


  (* keep_hierarchy = "yes" *) yshift
  yshift_27
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(yshift_27__ap_start),
    .ap_done(yshift_27__ap_done),
    .ap_idle(yshift_27__ap_idle),
    .ap_ready(yshift_27__ap_ready),
    .n(yshift_27___n__q0),
    .a_s_dout(qr27_vadd_bw__dout),
    .a_peek_dout(qr27_vadd_bw__dout),
    .a_s_empty_n(qr27_vadd_bw__empty_n),
    .a_peek_empty_n(qr27_vadd_bw__empty_n),
    .a_s_read(qr27_vadd_bw__read),
    .a_peek_read(),
    .b_din(qw27_vadd_bw__din),
    .b_full_n(qw27_vadd_bw__full_n),
    .b_write(qw27_vadd_bw__write)
  );


  (* keep_hierarchy = "yes" *) vadd_bw_fsm
  __tapa_fsm_unit
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(ap_start),
    .ap_done(ap_done),
    .ap_idle(ap_idle),
    .ap_ready(ap_ready),
    .n(n),
    .rmem0(rmem0),
    .rmem1(rmem1),
    .rmem2(rmem2),
    .rmem3(rmem3),
    .rmem4(rmem4),
    .rmem5(rmem5),
    .rmem6(rmem6),
    .rmem7(rmem7),
    .rmem8(rmem8),
    .rmem9(rmem9),
    .rmem10(rmem10),
    .rmem11(rmem11),
    .rmem12(rmem12),
    .rmem13(rmem13),
    .rmem14(rmem14),
    .rmem15(rmem15),
    .rmem16(rmem16),
    .rmem17(rmem17),
    .rmem18(rmem18),
    .rmem19(rmem19),
    .rmem20(rmem20),
    .rmem21(rmem21),
    .rmem22(rmem22),
    .rmem23(rmem23),
    .rmem24(rmem24),
    .rmem25(rmem25),
    .rmem26(rmem26),
    .rmem27(rmem27),
    .Mmap2Stream_0___n__q0(Mmap2Stream_0___n__q0),
    .Mmap2Stream_0___rmem0__q0(Mmap2Stream_0___rmem0__q0),
    .Mmap2Stream_0__ap_start(Mmap2Stream_0__ap_start),
    .Mmap2Stream_0__ap_ready(Mmap2Stream_0__ap_ready),
    .Mmap2Stream_0__ap_done(Mmap2Stream_0__ap_done),
    .Mmap2Stream_0__ap_idle(Mmap2Stream_0__ap_idle),
    .Mmap2Stream_1___n__q0(Mmap2Stream_1___n__q0),
    .Mmap2Stream_1___rmem1__q0(Mmap2Stream_1___rmem1__q0),
    .Mmap2Stream_1__ap_start(Mmap2Stream_1__ap_start),
    .Mmap2Stream_1__ap_ready(Mmap2Stream_1__ap_ready),
    .Mmap2Stream_1__ap_done(Mmap2Stream_1__ap_done),
    .Mmap2Stream_1__ap_idle(Mmap2Stream_1__ap_idle),
    .Mmap2Stream_2___n__q0(Mmap2Stream_2___n__q0),
    .Mmap2Stream_2___rmem2__q0(Mmap2Stream_2___rmem2__q0),
    .Mmap2Stream_2__ap_start(Mmap2Stream_2__ap_start),
    .Mmap2Stream_2__ap_ready(Mmap2Stream_2__ap_ready),
    .Mmap2Stream_2__ap_done(Mmap2Stream_2__ap_done),
    .Mmap2Stream_2__ap_idle(Mmap2Stream_2__ap_idle),
    .Mmap2Stream_3___n__q0(Mmap2Stream_3___n__q0),
    .Mmap2Stream_3___rmem3__q0(Mmap2Stream_3___rmem3__q0),
    .Mmap2Stream_3__ap_start(Mmap2Stream_3__ap_start),
    .Mmap2Stream_3__ap_ready(Mmap2Stream_3__ap_ready),
    .Mmap2Stream_3__ap_done(Mmap2Stream_3__ap_done),
    .Mmap2Stream_3__ap_idle(Mmap2Stream_3__ap_idle),
    .Mmap2Stream_4___n__q0(Mmap2Stream_4___n__q0),
    .Mmap2Stream_4___rmem4__q0(Mmap2Stream_4___rmem4__q0),
    .Mmap2Stream_4__ap_start(Mmap2Stream_4__ap_start),
    .Mmap2Stream_4__ap_ready(Mmap2Stream_4__ap_ready),
    .Mmap2Stream_4__ap_done(Mmap2Stream_4__ap_done),
    .Mmap2Stream_4__ap_idle(Mmap2Stream_4__ap_idle),
    .Mmap2Stream_5___n__q0(Mmap2Stream_5___n__q0),
    .Mmap2Stream_5___rmem5__q0(Mmap2Stream_5___rmem5__q0),
    .Mmap2Stream_5__ap_start(Mmap2Stream_5__ap_start),
    .Mmap2Stream_5__ap_ready(Mmap2Stream_5__ap_ready),
    .Mmap2Stream_5__ap_done(Mmap2Stream_5__ap_done),
    .Mmap2Stream_5__ap_idle(Mmap2Stream_5__ap_idle),
    .Mmap2Stream_6___n__q0(Mmap2Stream_6___n__q0),
    .Mmap2Stream_6___rmem6__q0(Mmap2Stream_6___rmem6__q0),
    .Mmap2Stream_6__ap_start(Mmap2Stream_6__ap_start),
    .Mmap2Stream_6__ap_ready(Mmap2Stream_6__ap_ready),
    .Mmap2Stream_6__ap_done(Mmap2Stream_6__ap_done),
    .Mmap2Stream_6__ap_idle(Mmap2Stream_6__ap_idle),
    .Mmap2Stream_7___n__q0(Mmap2Stream_7___n__q0),
    .Mmap2Stream_7___rmem7__q0(Mmap2Stream_7___rmem7__q0),
    .Mmap2Stream_7__ap_start(Mmap2Stream_7__ap_start),
    .Mmap2Stream_7__ap_ready(Mmap2Stream_7__ap_ready),
    .Mmap2Stream_7__ap_done(Mmap2Stream_7__ap_done),
    .Mmap2Stream_7__ap_idle(Mmap2Stream_7__ap_idle),
    .Mmap2Stream_8___n__q0(Mmap2Stream_8___n__q0),
    .Mmap2Stream_8___rmem8__q0(Mmap2Stream_8___rmem8__q0),
    .Mmap2Stream_8__ap_start(Mmap2Stream_8__ap_start),
    .Mmap2Stream_8__ap_ready(Mmap2Stream_8__ap_ready),
    .Mmap2Stream_8__ap_done(Mmap2Stream_8__ap_done),
    .Mmap2Stream_8__ap_idle(Mmap2Stream_8__ap_idle),
    .Mmap2Stream_9___n__q0(Mmap2Stream_9___n__q0),
    .Mmap2Stream_9___rmem9__q0(Mmap2Stream_9___rmem9__q0),
    .Mmap2Stream_9__ap_start(Mmap2Stream_9__ap_start),
    .Mmap2Stream_9__ap_ready(Mmap2Stream_9__ap_ready),
    .Mmap2Stream_9__ap_done(Mmap2Stream_9__ap_done),
    .Mmap2Stream_9__ap_idle(Mmap2Stream_9__ap_idle),
    .Mmap2Stream_10___n__q0(Mmap2Stream_10___n__q0),
    .Mmap2Stream_10___rmem10__q0(Mmap2Stream_10___rmem10__q0),
    .Mmap2Stream_10__ap_start(Mmap2Stream_10__ap_start),
    .Mmap2Stream_10__ap_ready(Mmap2Stream_10__ap_ready),
    .Mmap2Stream_10__ap_done(Mmap2Stream_10__ap_done),
    .Mmap2Stream_10__ap_idle(Mmap2Stream_10__ap_idle),
    .Mmap2Stream_11___n__q0(Mmap2Stream_11___n__q0),
    .Mmap2Stream_11___rmem11__q0(Mmap2Stream_11___rmem11__q0),
    .Mmap2Stream_11__ap_start(Mmap2Stream_11__ap_start),
    .Mmap2Stream_11__ap_ready(Mmap2Stream_11__ap_ready),
    .Mmap2Stream_11__ap_done(Mmap2Stream_11__ap_done),
    .Mmap2Stream_11__ap_idle(Mmap2Stream_11__ap_idle),
    .Mmap2Stream_12___n__q0(Mmap2Stream_12___n__q0),
    .Mmap2Stream_12___rmem12__q0(Mmap2Stream_12___rmem12__q0),
    .Mmap2Stream_12__ap_start(Mmap2Stream_12__ap_start),
    .Mmap2Stream_12__ap_ready(Mmap2Stream_12__ap_ready),
    .Mmap2Stream_12__ap_done(Mmap2Stream_12__ap_done),
    .Mmap2Stream_12__ap_idle(Mmap2Stream_12__ap_idle),
    .Mmap2Stream_13___n__q0(Mmap2Stream_13___n__q0),
    .Mmap2Stream_13___rmem13__q0(Mmap2Stream_13___rmem13__q0),
    .Mmap2Stream_13__ap_start(Mmap2Stream_13__ap_start),
    .Mmap2Stream_13__ap_ready(Mmap2Stream_13__ap_ready),
    .Mmap2Stream_13__ap_done(Mmap2Stream_13__ap_done),
    .Mmap2Stream_13__ap_idle(Mmap2Stream_13__ap_idle),
    .Mmap2Stream_14___n__q0(Mmap2Stream_14___n__q0),
    .Mmap2Stream_14___rmem14__q0(Mmap2Stream_14___rmem14__q0),
    .Mmap2Stream_14__ap_start(Mmap2Stream_14__ap_start),
    .Mmap2Stream_14__ap_ready(Mmap2Stream_14__ap_ready),
    .Mmap2Stream_14__ap_done(Mmap2Stream_14__ap_done),
    .Mmap2Stream_14__ap_idle(Mmap2Stream_14__ap_idle),
    .Mmap2Stream_15___n__q0(Mmap2Stream_15___n__q0),
    .Mmap2Stream_15___rmem15__q0(Mmap2Stream_15___rmem15__q0),
    .Mmap2Stream_15__ap_start(Mmap2Stream_15__ap_start),
    .Mmap2Stream_15__ap_ready(Mmap2Stream_15__ap_ready),
    .Mmap2Stream_15__ap_done(Mmap2Stream_15__ap_done),
    .Mmap2Stream_15__ap_idle(Mmap2Stream_15__ap_idle),
    .Mmap2Stream_16___n__q0(Mmap2Stream_16___n__q0),
    .Mmap2Stream_16___rmem16__q0(Mmap2Stream_16___rmem16__q0),
    .Mmap2Stream_16__ap_start(Mmap2Stream_16__ap_start),
    .Mmap2Stream_16__ap_ready(Mmap2Stream_16__ap_ready),
    .Mmap2Stream_16__ap_done(Mmap2Stream_16__ap_done),
    .Mmap2Stream_16__ap_idle(Mmap2Stream_16__ap_idle),
    .Mmap2Stream_17___n__q0(Mmap2Stream_17___n__q0),
    .Mmap2Stream_17___rmem17__q0(Mmap2Stream_17___rmem17__q0),
    .Mmap2Stream_17__ap_start(Mmap2Stream_17__ap_start),
    .Mmap2Stream_17__ap_ready(Mmap2Stream_17__ap_ready),
    .Mmap2Stream_17__ap_done(Mmap2Stream_17__ap_done),
    .Mmap2Stream_17__ap_idle(Mmap2Stream_17__ap_idle),
    .Mmap2Stream_18___n__q0(Mmap2Stream_18___n__q0),
    .Mmap2Stream_18___rmem18__q0(Mmap2Stream_18___rmem18__q0),
    .Mmap2Stream_18__ap_start(Mmap2Stream_18__ap_start),
    .Mmap2Stream_18__ap_ready(Mmap2Stream_18__ap_ready),
    .Mmap2Stream_18__ap_done(Mmap2Stream_18__ap_done),
    .Mmap2Stream_18__ap_idle(Mmap2Stream_18__ap_idle),
    .Mmap2Stream_19___n__q0(Mmap2Stream_19___n__q0),
    .Mmap2Stream_19___rmem19__q0(Mmap2Stream_19___rmem19__q0),
    .Mmap2Stream_19__ap_start(Mmap2Stream_19__ap_start),
    .Mmap2Stream_19__ap_ready(Mmap2Stream_19__ap_ready),
    .Mmap2Stream_19__ap_done(Mmap2Stream_19__ap_done),
    .Mmap2Stream_19__ap_idle(Mmap2Stream_19__ap_idle),
    .Mmap2Stream_20___n__q0(Mmap2Stream_20___n__q0),
    .Mmap2Stream_20___rmem20__q0(Mmap2Stream_20___rmem20__q0),
    .Mmap2Stream_20__ap_start(Mmap2Stream_20__ap_start),
    .Mmap2Stream_20__ap_ready(Mmap2Stream_20__ap_ready),
    .Mmap2Stream_20__ap_done(Mmap2Stream_20__ap_done),
    .Mmap2Stream_20__ap_idle(Mmap2Stream_20__ap_idle),
    .Mmap2Stream_21___n__q0(Mmap2Stream_21___n__q0),
    .Mmap2Stream_21___rmem21__q0(Mmap2Stream_21___rmem21__q0),
    .Mmap2Stream_21__ap_start(Mmap2Stream_21__ap_start),
    .Mmap2Stream_21__ap_ready(Mmap2Stream_21__ap_ready),
    .Mmap2Stream_21__ap_done(Mmap2Stream_21__ap_done),
    .Mmap2Stream_21__ap_idle(Mmap2Stream_21__ap_idle),
    .Mmap2Stream_22___n__q0(Mmap2Stream_22___n__q0),
    .Mmap2Stream_22___rmem22__q0(Mmap2Stream_22___rmem22__q0),
    .Mmap2Stream_22__ap_start(Mmap2Stream_22__ap_start),
    .Mmap2Stream_22__ap_ready(Mmap2Stream_22__ap_ready),
    .Mmap2Stream_22__ap_done(Mmap2Stream_22__ap_done),
    .Mmap2Stream_22__ap_idle(Mmap2Stream_22__ap_idle),
    .Mmap2Stream_23___n__q0(Mmap2Stream_23___n__q0),
    .Mmap2Stream_23___rmem23__q0(Mmap2Stream_23___rmem23__q0),
    .Mmap2Stream_23__ap_start(Mmap2Stream_23__ap_start),
    .Mmap2Stream_23__ap_ready(Mmap2Stream_23__ap_ready),
    .Mmap2Stream_23__ap_done(Mmap2Stream_23__ap_done),
    .Mmap2Stream_23__ap_idle(Mmap2Stream_23__ap_idle),
    .Mmap2Stream_24___n__q0(Mmap2Stream_24___n__q0),
    .Mmap2Stream_24___rmem24__q0(Mmap2Stream_24___rmem24__q0),
    .Mmap2Stream_24__ap_start(Mmap2Stream_24__ap_start),
    .Mmap2Stream_24__ap_ready(Mmap2Stream_24__ap_ready),
    .Mmap2Stream_24__ap_done(Mmap2Stream_24__ap_done),
    .Mmap2Stream_24__ap_idle(Mmap2Stream_24__ap_idle),
    .Mmap2Stream_25___n__q0(Mmap2Stream_25___n__q0),
    .Mmap2Stream_25___rmem25__q0(Mmap2Stream_25___rmem25__q0),
    .Mmap2Stream_25__ap_start(Mmap2Stream_25__ap_start),
    .Mmap2Stream_25__ap_ready(Mmap2Stream_25__ap_ready),
    .Mmap2Stream_25__ap_done(Mmap2Stream_25__ap_done),
    .Mmap2Stream_25__ap_idle(Mmap2Stream_25__ap_idle),
    .Mmap2Stream_26___n__q0(Mmap2Stream_26___n__q0),
    .Mmap2Stream_26___rmem26__q0(Mmap2Stream_26___rmem26__q0),
    .Mmap2Stream_26__ap_start(Mmap2Stream_26__ap_start),
    .Mmap2Stream_26__ap_ready(Mmap2Stream_26__ap_ready),
    .Mmap2Stream_26__ap_done(Mmap2Stream_26__ap_done),
    .Mmap2Stream_26__ap_idle(Mmap2Stream_26__ap_idle),
    .Mmap2Stream_27___n__q0(Mmap2Stream_27___n__q0),
    .Mmap2Stream_27___rmem27__q0(Mmap2Stream_27___rmem27__q0),
    .Mmap2Stream_27__ap_start(Mmap2Stream_27__ap_start),
    .Mmap2Stream_27__ap_ready(Mmap2Stream_27__ap_ready),
    .Mmap2Stream_27__ap_done(Mmap2Stream_27__ap_done),
    .Mmap2Stream_27__ap_idle(Mmap2Stream_27__ap_idle),
    .Stream2Mmap_0___n__q0(Stream2Mmap_0___n__q0),
    .Stream2Mmap_0___rmem0__q0(Stream2Mmap_0___rmem0__q0),
    .Stream2Mmap_0__ap_start(Stream2Mmap_0__ap_start),
    .Stream2Mmap_0__ap_ready(Stream2Mmap_0__ap_ready),
    .Stream2Mmap_0__ap_done(Stream2Mmap_0__ap_done),
    .Stream2Mmap_0__ap_idle(Stream2Mmap_0__ap_idle),
    .Stream2Mmap_1___n__q0(Stream2Mmap_1___n__q0),
    .Stream2Mmap_1___rmem1__q0(Stream2Mmap_1___rmem1__q0),
    .Stream2Mmap_1__ap_start(Stream2Mmap_1__ap_start),
    .Stream2Mmap_1__ap_ready(Stream2Mmap_1__ap_ready),
    .Stream2Mmap_1__ap_done(Stream2Mmap_1__ap_done),
    .Stream2Mmap_1__ap_idle(Stream2Mmap_1__ap_idle),
    .Stream2Mmap_2___n__q0(Stream2Mmap_2___n__q0),
    .Stream2Mmap_2___rmem2__q0(Stream2Mmap_2___rmem2__q0),
    .Stream2Mmap_2__ap_start(Stream2Mmap_2__ap_start),
    .Stream2Mmap_2__ap_ready(Stream2Mmap_2__ap_ready),
    .Stream2Mmap_2__ap_done(Stream2Mmap_2__ap_done),
    .Stream2Mmap_2__ap_idle(Stream2Mmap_2__ap_idle),
    .Stream2Mmap_3___n__q0(Stream2Mmap_3___n__q0),
    .Stream2Mmap_3___rmem3__q0(Stream2Mmap_3___rmem3__q0),
    .Stream2Mmap_3__ap_start(Stream2Mmap_3__ap_start),
    .Stream2Mmap_3__ap_ready(Stream2Mmap_3__ap_ready),
    .Stream2Mmap_3__ap_done(Stream2Mmap_3__ap_done),
    .Stream2Mmap_3__ap_idle(Stream2Mmap_3__ap_idle),
    .Stream2Mmap_4___n__q0(Stream2Mmap_4___n__q0),
    .Stream2Mmap_4___rmem4__q0(Stream2Mmap_4___rmem4__q0),
    .Stream2Mmap_4__ap_start(Stream2Mmap_4__ap_start),
    .Stream2Mmap_4__ap_ready(Stream2Mmap_4__ap_ready),
    .Stream2Mmap_4__ap_done(Stream2Mmap_4__ap_done),
    .Stream2Mmap_4__ap_idle(Stream2Mmap_4__ap_idle),
    .Stream2Mmap_5___n__q0(Stream2Mmap_5___n__q0),
    .Stream2Mmap_5___rmem5__q0(Stream2Mmap_5___rmem5__q0),
    .Stream2Mmap_5__ap_start(Stream2Mmap_5__ap_start),
    .Stream2Mmap_5__ap_ready(Stream2Mmap_5__ap_ready),
    .Stream2Mmap_5__ap_done(Stream2Mmap_5__ap_done),
    .Stream2Mmap_5__ap_idle(Stream2Mmap_5__ap_idle),
    .Stream2Mmap_6___n__q0(Stream2Mmap_6___n__q0),
    .Stream2Mmap_6___rmem6__q0(Stream2Mmap_6___rmem6__q0),
    .Stream2Mmap_6__ap_start(Stream2Mmap_6__ap_start),
    .Stream2Mmap_6__ap_ready(Stream2Mmap_6__ap_ready),
    .Stream2Mmap_6__ap_done(Stream2Mmap_6__ap_done),
    .Stream2Mmap_6__ap_idle(Stream2Mmap_6__ap_idle),
    .Stream2Mmap_7___n__q0(Stream2Mmap_7___n__q0),
    .Stream2Mmap_7___rmem7__q0(Stream2Mmap_7___rmem7__q0),
    .Stream2Mmap_7__ap_start(Stream2Mmap_7__ap_start),
    .Stream2Mmap_7__ap_ready(Stream2Mmap_7__ap_ready),
    .Stream2Mmap_7__ap_done(Stream2Mmap_7__ap_done),
    .Stream2Mmap_7__ap_idle(Stream2Mmap_7__ap_idle),
    .Stream2Mmap_8___n__q0(Stream2Mmap_8___n__q0),
    .Stream2Mmap_8___rmem8__q0(Stream2Mmap_8___rmem8__q0),
    .Stream2Mmap_8__ap_start(Stream2Mmap_8__ap_start),
    .Stream2Mmap_8__ap_ready(Stream2Mmap_8__ap_ready),
    .Stream2Mmap_8__ap_done(Stream2Mmap_8__ap_done),
    .Stream2Mmap_8__ap_idle(Stream2Mmap_8__ap_idle),
    .Stream2Mmap_9___n__q0(Stream2Mmap_9___n__q0),
    .Stream2Mmap_9___rmem9__q0(Stream2Mmap_9___rmem9__q0),
    .Stream2Mmap_9__ap_start(Stream2Mmap_9__ap_start),
    .Stream2Mmap_9__ap_ready(Stream2Mmap_9__ap_ready),
    .Stream2Mmap_9__ap_done(Stream2Mmap_9__ap_done),
    .Stream2Mmap_9__ap_idle(Stream2Mmap_9__ap_idle),
    .Stream2Mmap_10___n__q0(Stream2Mmap_10___n__q0),
    .Stream2Mmap_10___rmem10__q0(Stream2Mmap_10___rmem10__q0),
    .Stream2Mmap_10__ap_start(Stream2Mmap_10__ap_start),
    .Stream2Mmap_10__ap_ready(Stream2Mmap_10__ap_ready),
    .Stream2Mmap_10__ap_done(Stream2Mmap_10__ap_done),
    .Stream2Mmap_10__ap_idle(Stream2Mmap_10__ap_idle),
    .Stream2Mmap_11___n__q0(Stream2Mmap_11___n__q0),
    .Stream2Mmap_11___rmem11__q0(Stream2Mmap_11___rmem11__q0),
    .Stream2Mmap_11__ap_start(Stream2Mmap_11__ap_start),
    .Stream2Mmap_11__ap_ready(Stream2Mmap_11__ap_ready),
    .Stream2Mmap_11__ap_done(Stream2Mmap_11__ap_done),
    .Stream2Mmap_11__ap_idle(Stream2Mmap_11__ap_idle),
    .Stream2Mmap_12___n__q0(Stream2Mmap_12___n__q0),
    .Stream2Mmap_12___rmem12__q0(Stream2Mmap_12___rmem12__q0),
    .Stream2Mmap_12__ap_start(Stream2Mmap_12__ap_start),
    .Stream2Mmap_12__ap_ready(Stream2Mmap_12__ap_ready),
    .Stream2Mmap_12__ap_done(Stream2Mmap_12__ap_done),
    .Stream2Mmap_12__ap_idle(Stream2Mmap_12__ap_idle),
    .Stream2Mmap_13___n__q0(Stream2Mmap_13___n__q0),
    .Stream2Mmap_13___rmem13__q0(Stream2Mmap_13___rmem13__q0),
    .Stream2Mmap_13__ap_start(Stream2Mmap_13__ap_start),
    .Stream2Mmap_13__ap_ready(Stream2Mmap_13__ap_ready),
    .Stream2Mmap_13__ap_done(Stream2Mmap_13__ap_done),
    .Stream2Mmap_13__ap_idle(Stream2Mmap_13__ap_idle),
    .Stream2Mmap_14___n__q0(Stream2Mmap_14___n__q0),
    .Stream2Mmap_14___rmem14__q0(Stream2Mmap_14___rmem14__q0),
    .Stream2Mmap_14__ap_start(Stream2Mmap_14__ap_start),
    .Stream2Mmap_14__ap_ready(Stream2Mmap_14__ap_ready),
    .Stream2Mmap_14__ap_done(Stream2Mmap_14__ap_done),
    .Stream2Mmap_14__ap_idle(Stream2Mmap_14__ap_idle),
    .Stream2Mmap_15___n__q0(Stream2Mmap_15___n__q0),
    .Stream2Mmap_15___rmem15__q0(Stream2Mmap_15___rmem15__q0),
    .Stream2Mmap_15__ap_start(Stream2Mmap_15__ap_start),
    .Stream2Mmap_15__ap_ready(Stream2Mmap_15__ap_ready),
    .Stream2Mmap_15__ap_done(Stream2Mmap_15__ap_done),
    .Stream2Mmap_15__ap_idle(Stream2Mmap_15__ap_idle),
    .Stream2Mmap_16___n__q0(Stream2Mmap_16___n__q0),
    .Stream2Mmap_16___rmem16__q0(Stream2Mmap_16___rmem16__q0),
    .Stream2Mmap_16__ap_start(Stream2Mmap_16__ap_start),
    .Stream2Mmap_16__ap_ready(Stream2Mmap_16__ap_ready),
    .Stream2Mmap_16__ap_done(Stream2Mmap_16__ap_done),
    .Stream2Mmap_16__ap_idle(Stream2Mmap_16__ap_idle),
    .Stream2Mmap_17___n__q0(Stream2Mmap_17___n__q0),
    .Stream2Mmap_17___rmem17__q0(Stream2Mmap_17___rmem17__q0),
    .Stream2Mmap_17__ap_start(Stream2Mmap_17__ap_start),
    .Stream2Mmap_17__ap_ready(Stream2Mmap_17__ap_ready),
    .Stream2Mmap_17__ap_done(Stream2Mmap_17__ap_done),
    .Stream2Mmap_17__ap_idle(Stream2Mmap_17__ap_idle),
    .Stream2Mmap_18___n__q0(Stream2Mmap_18___n__q0),
    .Stream2Mmap_18___rmem18__q0(Stream2Mmap_18___rmem18__q0),
    .Stream2Mmap_18__ap_start(Stream2Mmap_18__ap_start),
    .Stream2Mmap_18__ap_ready(Stream2Mmap_18__ap_ready),
    .Stream2Mmap_18__ap_done(Stream2Mmap_18__ap_done),
    .Stream2Mmap_18__ap_idle(Stream2Mmap_18__ap_idle),
    .Stream2Mmap_19___n__q0(Stream2Mmap_19___n__q0),
    .Stream2Mmap_19___rmem19__q0(Stream2Mmap_19___rmem19__q0),
    .Stream2Mmap_19__ap_start(Stream2Mmap_19__ap_start),
    .Stream2Mmap_19__ap_ready(Stream2Mmap_19__ap_ready),
    .Stream2Mmap_19__ap_done(Stream2Mmap_19__ap_done),
    .Stream2Mmap_19__ap_idle(Stream2Mmap_19__ap_idle),
    .Stream2Mmap_20___n__q0(Stream2Mmap_20___n__q0),
    .Stream2Mmap_20___rmem20__q0(Stream2Mmap_20___rmem20__q0),
    .Stream2Mmap_20__ap_start(Stream2Mmap_20__ap_start),
    .Stream2Mmap_20__ap_ready(Stream2Mmap_20__ap_ready),
    .Stream2Mmap_20__ap_done(Stream2Mmap_20__ap_done),
    .Stream2Mmap_20__ap_idle(Stream2Mmap_20__ap_idle),
    .Stream2Mmap_21___n__q0(Stream2Mmap_21___n__q0),
    .Stream2Mmap_21___rmem21__q0(Stream2Mmap_21___rmem21__q0),
    .Stream2Mmap_21__ap_start(Stream2Mmap_21__ap_start),
    .Stream2Mmap_21__ap_ready(Stream2Mmap_21__ap_ready),
    .Stream2Mmap_21__ap_done(Stream2Mmap_21__ap_done),
    .Stream2Mmap_21__ap_idle(Stream2Mmap_21__ap_idle),
    .Stream2Mmap_22___n__q0(Stream2Mmap_22___n__q0),
    .Stream2Mmap_22___rmem22__q0(Stream2Mmap_22___rmem22__q0),
    .Stream2Mmap_22__ap_start(Stream2Mmap_22__ap_start),
    .Stream2Mmap_22__ap_ready(Stream2Mmap_22__ap_ready),
    .Stream2Mmap_22__ap_done(Stream2Mmap_22__ap_done),
    .Stream2Mmap_22__ap_idle(Stream2Mmap_22__ap_idle),
    .Stream2Mmap_23___n__q0(Stream2Mmap_23___n__q0),
    .Stream2Mmap_23___rmem23__q0(Stream2Mmap_23___rmem23__q0),
    .Stream2Mmap_23__ap_start(Stream2Mmap_23__ap_start),
    .Stream2Mmap_23__ap_ready(Stream2Mmap_23__ap_ready),
    .Stream2Mmap_23__ap_done(Stream2Mmap_23__ap_done),
    .Stream2Mmap_23__ap_idle(Stream2Mmap_23__ap_idle),
    .Stream2Mmap_24___n__q0(Stream2Mmap_24___n__q0),
    .Stream2Mmap_24___rmem24__q0(Stream2Mmap_24___rmem24__q0),
    .Stream2Mmap_24__ap_start(Stream2Mmap_24__ap_start),
    .Stream2Mmap_24__ap_ready(Stream2Mmap_24__ap_ready),
    .Stream2Mmap_24__ap_done(Stream2Mmap_24__ap_done),
    .Stream2Mmap_24__ap_idle(Stream2Mmap_24__ap_idle),
    .Stream2Mmap_25___n__q0(Stream2Mmap_25___n__q0),
    .Stream2Mmap_25___rmem25__q0(Stream2Mmap_25___rmem25__q0),
    .Stream2Mmap_25__ap_start(Stream2Mmap_25__ap_start),
    .Stream2Mmap_25__ap_ready(Stream2Mmap_25__ap_ready),
    .Stream2Mmap_25__ap_done(Stream2Mmap_25__ap_done),
    .Stream2Mmap_25__ap_idle(Stream2Mmap_25__ap_idle),
    .Stream2Mmap_26___n__q0(Stream2Mmap_26___n__q0),
    .Stream2Mmap_26___rmem26__q0(Stream2Mmap_26___rmem26__q0),
    .Stream2Mmap_26__ap_start(Stream2Mmap_26__ap_start),
    .Stream2Mmap_26__ap_ready(Stream2Mmap_26__ap_ready),
    .Stream2Mmap_26__ap_done(Stream2Mmap_26__ap_done),
    .Stream2Mmap_26__ap_idle(Stream2Mmap_26__ap_idle),
    .Stream2Mmap_27___n__q0(Stream2Mmap_27___n__q0),
    .Stream2Mmap_27___rmem27__q0(Stream2Mmap_27___rmem27__q0),
    .Stream2Mmap_27__ap_start(Stream2Mmap_27__ap_start),
    .Stream2Mmap_27__ap_ready(Stream2Mmap_27__ap_ready),
    .Stream2Mmap_27__ap_done(Stream2Mmap_27__ap_done),
    .Stream2Mmap_27__ap_idle(Stream2Mmap_27__ap_idle),
    .yshift_0___n__q0(yshift_0___n__q0),
    .yshift_0__ap_start(yshift_0__ap_start),
    .yshift_0__ap_ready(yshift_0__ap_ready),
    .yshift_0__ap_done(yshift_0__ap_done),
    .yshift_0__ap_idle(yshift_0__ap_idle),
    .yshift_1___n__q0(yshift_1___n__q0),
    .yshift_1__ap_start(yshift_1__ap_start),
    .yshift_1__ap_ready(yshift_1__ap_ready),
    .yshift_1__ap_done(yshift_1__ap_done),
    .yshift_1__ap_idle(yshift_1__ap_idle),
    .yshift_2___n__q0(yshift_2___n__q0),
    .yshift_2__ap_start(yshift_2__ap_start),
    .yshift_2__ap_ready(yshift_2__ap_ready),
    .yshift_2__ap_done(yshift_2__ap_done),
    .yshift_2__ap_idle(yshift_2__ap_idle),
    .yshift_3___n__q0(yshift_3___n__q0),
    .yshift_3__ap_start(yshift_3__ap_start),
    .yshift_3__ap_ready(yshift_3__ap_ready),
    .yshift_3__ap_done(yshift_3__ap_done),
    .yshift_3__ap_idle(yshift_3__ap_idle),
    .yshift_4___n__q0(yshift_4___n__q0),
    .yshift_4__ap_start(yshift_4__ap_start),
    .yshift_4__ap_ready(yshift_4__ap_ready),
    .yshift_4__ap_done(yshift_4__ap_done),
    .yshift_4__ap_idle(yshift_4__ap_idle),
    .yshift_5___n__q0(yshift_5___n__q0),
    .yshift_5__ap_start(yshift_5__ap_start),
    .yshift_5__ap_ready(yshift_5__ap_ready),
    .yshift_5__ap_done(yshift_5__ap_done),
    .yshift_5__ap_idle(yshift_5__ap_idle),
    .yshift_6___n__q0(yshift_6___n__q0),
    .yshift_6__ap_start(yshift_6__ap_start),
    .yshift_6__ap_ready(yshift_6__ap_ready),
    .yshift_6__ap_done(yshift_6__ap_done),
    .yshift_6__ap_idle(yshift_6__ap_idle),
    .yshift_7___n__q0(yshift_7___n__q0),
    .yshift_7__ap_start(yshift_7__ap_start),
    .yshift_7__ap_ready(yshift_7__ap_ready),
    .yshift_7__ap_done(yshift_7__ap_done),
    .yshift_7__ap_idle(yshift_7__ap_idle),
    .yshift_8___n__q0(yshift_8___n__q0),
    .yshift_8__ap_start(yshift_8__ap_start),
    .yshift_8__ap_ready(yshift_8__ap_ready),
    .yshift_8__ap_done(yshift_8__ap_done),
    .yshift_8__ap_idle(yshift_8__ap_idle),
    .yshift_9___n__q0(yshift_9___n__q0),
    .yshift_9__ap_start(yshift_9__ap_start),
    .yshift_9__ap_ready(yshift_9__ap_ready),
    .yshift_9__ap_done(yshift_9__ap_done),
    .yshift_9__ap_idle(yshift_9__ap_idle),
    .yshift_10___n__q0(yshift_10___n__q0),
    .yshift_10__ap_start(yshift_10__ap_start),
    .yshift_10__ap_ready(yshift_10__ap_ready),
    .yshift_10__ap_done(yshift_10__ap_done),
    .yshift_10__ap_idle(yshift_10__ap_idle),
    .yshift_11___n__q0(yshift_11___n__q0),
    .yshift_11__ap_start(yshift_11__ap_start),
    .yshift_11__ap_ready(yshift_11__ap_ready),
    .yshift_11__ap_done(yshift_11__ap_done),
    .yshift_11__ap_idle(yshift_11__ap_idle),
    .yshift_12___n__q0(yshift_12___n__q0),
    .yshift_12__ap_start(yshift_12__ap_start),
    .yshift_12__ap_ready(yshift_12__ap_ready),
    .yshift_12__ap_done(yshift_12__ap_done),
    .yshift_12__ap_idle(yshift_12__ap_idle),
    .yshift_13___n__q0(yshift_13___n__q0),
    .yshift_13__ap_start(yshift_13__ap_start),
    .yshift_13__ap_ready(yshift_13__ap_ready),
    .yshift_13__ap_done(yshift_13__ap_done),
    .yshift_13__ap_idle(yshift_13__ap_idle),
    .yshift_14___n__q0(yshift_14___n__q0),
    .yshift_14__ap_start(yshift_14__ap_start),
    .yshift_14__ap_ready(yshift_14__ap_ready),
    .yshift_14__ap_done(yshift_14__ap_done),
    .yshift_14__ap_idle(yshift_14__ap_idle),
    .yshift_15___n__q0(yshift_15___n__q0),
    .yshift_15__ap_start(yshift_15__ap_start),
    .yshift_15__ap_ready(yshift_15__ap_ready),
    .yshift_15__ap_done(yshift_15__ap_done),
    .yshift_15__ap_idle(yshift_15__ap_idle),
    .yshift_16___n__q0(yshift_16___n__q0),
    .yshift_16__ap_start(yshift_16__ap_start),
    .yshift_16__ap_ready(yshift_16__ap_ready),
    .yshift_16__ap_done(yshift_16__ap_done),
    .yshift_16__ap_idle(yshift_16__ap_idle),
    .yshift_17___n__q0(yshift_17___n__q0),
    .yshift_17__ap_start(yshift_17__ap_start),
    .yshift_17__ap_ready(yshift_17__ap_ready),
    .yshift_17__ap_done(yshift_17__ap_done),
    .yshift_17__ap_idle(yshift_17__ap_idle),
    .yshift_18___n__q0(yshift_18___n__q0),
    .yshift_18__ap_start(yshift_18__ap_start),
    .yshift_18__ap_ready(yshift_18__ap_ready),
    .yshift_18__ap_done(yshift_18__ap_done),
    .yshift_18__ap_idle(yshift_18__ap_idle),
    .yshift_19___n__q0(yshift_19___n__q0),
    .yshift_19__ap_start(yshift_19__ap_start),
    .yshift_19__ap_ready(yshift_19__ap_ready),
    .yshift_19__ap_done(yshift_19__ap_done),
    .yshift_19__ap_idle(yshift_19__ap_idle),
    .yshift_20___n__q0(yshift_20___n__q0),
    .yshift_20__ap_start(yshift_20__ap_start),
    .yshift_20__ap_ready(yshift_20__ap_ready),
    .yshift_20__ap_done(yshift_20__ap_done),
    .yshift_20__ap_idle(yshift_20__ap_idle),
    .yshift_21___n__q0(yshift_21___n__q0),
    .yshift_21__ap_start(yshift_21__ap_start),
    .yshift_21__ap_ready(yshift_21__ap_ready),
    .yshift_21__ap_done(yshift_21__ap_done),
    .yshift_21__ap_idle(yshift_21__ap_idle),
    .yshift_22___n__q0(yshift_22___n__q0),
    .yshift_22__ap_start(yshift_22__ap_start),
    .yshift_22__ap_ready(yshift_22__ap_ready),
    .yshift_22__ap_done(yshift_22__ap_done),
    .yshift_22__ap_idle(yshift_22__ap_idle),
    .yshift_23___n__q0(yshift_23___n__q0),
    .yshift_23__ap_start(yshift_23__ap_start),
    .yshift_23__ap_ready(yshift_23__ap_ready),
    .yshift_23__ap_done(yshift_23__ap_done),
    .yshift_23__ap_idle(yshift_23__ap_idle),
    .yshift_24___n__q0(yshift_24___n__q0),
    .yshift_24__ap_start(yshift_24__ap_start),
    .yshift_24__ap_ready(yshift_24__ap_ready),
    .yshift_24__ap_done(yshift_24__ap_done),
    .yshift_24__ap_idle(yshift_24__ap_idle),
    .yshift_25___n__q0(yshift_25___n__q0),
    .yshift_25__ap_start(yshift_25__ap_start),
    .yshift_25__ap_ready(yshift_25__ap_ready),
    .yshift_25__ap_done(yshift_25__ap_done),
    .yshift_25__ap_idle(yshift_25__ap_idle),
    .yshift_26___n__q0(yshift_26___n__q0),
    .yshift_26__ap_start(yshift_26__ap_start),
    .yshift_26__ap_ready(yshift_26__ap_ready),
    .yshift_26__ap_done(yshift_26__ap_done),
    .yshift_26__ap_idle(yshift_26__ap_idle),
    .yshift_27___n__q0(yshift_27___n__q0),
    .yshift_27__ap_start(yshift_27__ap_start),
    .yshift_27__ap_ready(yshift_27__ap_ready),
    .yshift_27__ap_done(yshift_27__ap_done),
    .yshift_27__ap_idle(yshift_27__ap_idle)
  );

  assign ap_rst_n_inv = (~ap_rst_n);

endmodule
