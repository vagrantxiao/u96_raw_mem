

module vadd_bw_fsm
(
  ap_clk,
  ap_rst_n,
  ap_start,
  ap_ready,
  ap_done,
  ap_idle,
  n,
  rmem0,
  rmem1,
  rmem2,
  rmem3,
  rmem4,
  rmem5,
  rmem6,
  rmem7,
  rmem8,
  rmem9,
  rmem10,
  rmem11,
  rmem12,
  rmem13,
  rmem14,
  rmem15,
  rmem16,
  rmem17,
  rmem18,
  rmem19,
  rmem20,
  rmem21,
  rmem22,
  rmem23,
  rmem24,
  rmem25,
  rmem26,
  Mmap2Stream_0___n__q0,
  Mmap2Stream_0___rmem0__q0,
  Mmap2Stream_0__ap_start,
  Mmap2Stream_0__ap_ready,
  Mmap2Stream_0__ap_done,
  Mmap2Stream_0__ap_idle,
  Mmap2Stream_1___n__q0,
  Mmap2Stream_1___rmem1__q0,
  Mmap2Stream_1__ap_start,
  Mmap2Stream_1__ap_ready,
  Mmap2Stream_1__ap_done,
  Mmap2Stream_1__ap_idle,
  Mmap2Stream_2___n__q0,
  Mmap2Stream_2___rmem2__q0,
  Mmap2Stream_2__ap_start,
  Mmap2Stream_2__ap_ready,
  Mmap2Stream_2__ap_done,
  Mmap2Stream_2__ap_idle,
  Mmap2Stream_3___n__q0,
  Mmap2Stream_3___rmem3__q0,
  Mmap2Stream_3__ap_start,
  Mmap2Stream_3__ap_ready,
  Mmap2Stream_3__ap_done,
  Mmap2Stream_3__ap_idle,
  Mmap2Stream_4___n__q0,
  Mmap2Stream_4___rmem4__q0,
  Mmap2Stream_4__ap_start,
  Mmap2Stream_4__ap_ready,
  Mmap2Stream_4__ap_done,
  Mmap2Stream_4__ap_idle,
  Mmap2Stream_5___n__q0,
  Mmap2Stream_5___rmem5__q0,
  Mmap2Stream_5__ap_start,
  Mmap2Stream_5__ap_ready,
  Mmap2Stream_5__ap_done,
  Mmap2Stream_5__ap_idle,
  Mmap2Stream_6___n__q0,
  Mmap2Stream_6___rmem6__q0,
  Mmap2Stream_6__ap_start,
  Mmap2Stream_6__ap_ready,
  Mmap2Stream_6__ap_done,
  Mmap2Stream_6__ap_idle,
  Mmap2Stream_7___n__q0,
  Mmap2Stream_7___rmem7__q0,
  Mmap2Stream_7__ap_start,
  Mmap2Stream_7__ap_ready,
  Mmap2Stream_7__ap_done,
  Mmap2Stream_7__ap_idle,
  Mmap2Stream_8___n__q0,
  Mmap2Stream_8___rmem8__q0,
  Mmap2Stream_8__ap_start,
  Mmap2Stream_8__ap_ready,
  Mmap2Stream_8__ap_done,
  Mmap2Stream_8__ap_idle,
  Mmap2Stream_9___n__q0,
  Mmap2Stream_9___rmem9__q0,
  Mmap2Stream_9__ap_start,
  Mmap2Stream_9__ap_ready,
  Mmap2Stream_9__ap_done,
  Mmap2Stream_9__ap_idle,
  Mmap2Stream_10___n__q0,
  Mmap2Stream_10___rmem10__q0,
  Mmap2Stream_10__ap_start,
  Mmap2Stream_10__ap_ready,
  Mmap2Stream_10__ap_done,
  Mmap2Stream_10__ap_idle,
  Mmap2Stream_11___n__q0,
  Mmap2Stream_11___rmem11__q0,
  Mmap2Stream_11__ap_start,
  Mmap2Stream_11__ap_ready,
  Mmap2Stream_11__ap_done,
  Mmap2Stream_11__ap_idle,
  Mmap2Stream_12___n__q0,
  Mmap2Stream_12___rmem12__q0,
  Mmap2Stream_12__ap_start,
  Mmap2Stream_12__ap_ready,
  Mmap2Stream_12__ap_done,
  Mmap2Stream_12__ap_idle,
  Mmap2Stream_13___n__q0,
  Mmap2Stream_13___rmem13__q0,
  Mmap2Stream_13__ap_start,
  Mmap2Stream_13__ap_ready,
  Mmap2Stream_13__ap_done,
  Mmap2Stream_13__ap_idle,
  Mmap2Stream_14___n__q0,
  Mmap2Stream_14___rmem14__q0,
  Mmap2Stream_14__ap_start,
  Mmap2Stream_14__ap_ready,
  Mmap2Stream_14__ap_done,
  Mmap2Stream_14__ap_idle,
  Mmap2Stream_15___n__q0,
  Mmap2Stream_15___rmem15__q0,
  Mmap2Stream_15__ap_start,
  Mmap2Stream_15__ap_ready,
  Mmap2Stream_15__ap_done,
  Mmap2Stream_15__ap_idle,
  Mmap2Stream_16___n__q0,
  Mmap2Stream_16___rmem16__q0,
  Mmap2Stream_16__ap_start,
  Mmap2Stream_16__ap_ready,
  Mmap2Stream_16__ap_done,
  Mmap2Stream_16__ap_idle,
  Mmap2Stream_17___n__q0,
  Mmap2Stream_17___rmem17__q0,
  Mmap2Stream_17__ap_start,
  Mmap2Stream_17__ap_ready,
  Mmap2Stream_17__ap_done,
  Mmap2Stream_17__ap_idle,
  Mmap2Stream_18___n__q0,
  Mmap2Stream_18___rmem18__q0,
  Mmap2Stream_18__ap_start,
  Mmap2Stream_18__ap_ready,
  Mmap2Stream_18__ap_done,
  Mmap2Stream_18__ap_idle,
  Mmap2Stream_19___n__q0,
  Mmap2Stream_19___rmem19__q0,
  Mmap2Stream_19__ap_start,
  Mmap2Stream_19__ap_ready,
  Mmap2Stream_19__ap_done,
  Mmap2Stream_19__ap_idle,
  Mmap2Stream_20___n__q0,
  Mmap2Stream_20___rmem20__q0,
  Mmap2Stream_20__ap_start,
  Mmap2Stream_20__ap_ready,
  Mmap2Stream_20__ap_done,
  Mmap2Stream_20__ap_idle,
  Mmap2Stream_21___n__q0,
  Mmap2Stream_21___rmem21__q0,
  Mmap2Stream_21__ap_start,
  Mmap2Stream_21__ap_ready,
  Mmap2Stream_21__ap_done,
  Mmap2Stream_21__ap_idle,
  Mmap2Stream_22___n__q0,
  Mmap2Stream_22___rmem22__q0,
  Mmap2Stream_22__ap_start,
  Mmap2Stream_22__ap_ready,
  Mmap2Stream_22__ap_done,
  Mmap2Stream_22__ap_idle,
  Mmap2Stream_23___n__q0,
  Mmap2Stream_23___rmem23__q0,
  Mmap2Stream_23__ap_start,
  Mmap2Stream_23__ap_ready,
  Mmap2Stream_23__ap_done,
  Mmap2Stream_23__ap_idle,
  Mmap2Stream_24___n__q0,
  Mmap2Stream_24___rmem24__q0,
  Mmap2Stream_24__ap_start,
  Mmap2Stream_24__ap_ready,
  Mmap2Stream_24__ap_done,
  Mmap2Stream_24__ap_idle,
  Mmap2Stream_25___n__q0,
  Mmap2Stream_25___rmem25__q0,
  Mmap2Stream_25__ap_start,
  Mmap2Stream_25__ap_ready,
  Mmap2Stream_25__ap_done,
  Mmap2Stream_25__ap_idle,
  Mmap2Stream_26___n__q0,
  Mmap2Stream_26___rmem26__q0,
  Mmap2Stream_26__ap_start,
  Mmap2Stream_26__ap_ready,
  Mmap2Stream_26__ap_done,
  Mmap2Stream_26__ap_idle,
  Stream2Mmap_0___n__q0,
  Stream2Mmap_0___rmem0__q0,
  Stream2Mmap_0__ap_start,
  Stream2Mmap_0__ap_ready,
  Stream2Mmap_0__ap_done,
  Stream2Mmap_0__ap_idle,
  Stream2Mmap_1___n__q0,
  Stream2Mmap_1___rmem1__q0,
  Stream2Mmap_1__ap_start,
  Stream2Mmap_1__ap_ready,
  Stream2Mmap_1__ap_done,
  Stream2Mmap_1__ap_idle,
  Stream2Mmap_2___n__q0,
  Stream2Mmap_2___rmem2__q0,
  Stream2Mmap_2__ap_start,
  Stream2Mmap_2__ap_ready,
  Stream2Mmap_2__ap_done,
  Stream2Mmap_2__ap_idle,
  Stream2Mmap_3___n__q0,
  Stream2Mmap_3___rmem3__q0,
  Stream2Mmap_3__ap_start,
  Stream2Mmap_3__ap_ready,
  Stream2Mmap_3__ap_done,
  Stream2Mmap_3__ap_idle,
  Stream2Mmap_4___n__q0,
  Stream2Mmap_4___rmem4__q0,
  Stream2Mmap_4__ap_start,
  Stream2Mmap_4__ap_ready,
  Stream2Mmap_4__ap_done,
  Stream2Mmap_4__ap_idle,
  Stream2Mmap_5___n__q0,
  Stream2Mmap_5___rmem5__q0,
  Stream2Mmap_5__ap_start,
  Stream2Mmap_5__ap_ready,
  Stream2Mmap_5__ap_done,
  Stream2Mmap_5__ap_idle,
  Stream2Mmap_6___n__q0,
  Stream2Mmap_6___rmem6__q0,
  Stream2Mmap_6__ap_start,
  Stream2Mmap_6__ap_ready,
  Stream2Mmap_6__ap_done,
  Stream2Mmap_6__ap_idle,
  Stream2Mmap_7___n__q0,
  Stream2Mmap_7___rmem7__q0,
  Stream2Mmap_7__ap_start,
  Stream2Mmap_7__ap_ready,
  Stream2Mmap_7__ap_done,
  Stream2Mmap_7__ap_idle,
  Stream2Mmap_8___n__q0,
  Stream2Mmap_8___rmem8__q0,
  Stream2Mmap_8__ap_start,
  Stream2Mmap_8__ap_ready,
  Stream2Mmap_8__ap_done,
  Stream2Mmap_8__ap_idle,
  Stream2Mmap_9___n__q0,
  Stream2Mmap_9___rmem9__q0,
  Stream2Mmap_9__ap_start,
  Stream2Mmap_9__ap_ready,
  Stream2Mmap_9__ap_done,
  Stream2Mmap_9__ap_idle,
  Stream2Mmap_10___n__q0,
  Stream2Mmap_10___rmem10__q0,
  Stream2Mmap_10__ap_start,
  Stream2Mmap_10__ap_ready,
  Stream2Mmap_10__ap_done,
  Stream2Mmap_10__ap_idle,
  Stream2Mmap_11___n__q0,
  Stream2Mmap_11___rmem11__q0,
  Stream2Mmap_11__ap_start,
  Stream2Mmap_11__ap_ready,
  Stream2Mmap_11__ap_done,
  Stream2Mmap_11__ap_idle,
  Stream2Mmap_12___n__q0,
  Stream2Mmap_12___rmem12__q0,
  Stream2Mmap_12__ap_start,
  Stream2Mmap_12__ap_ready,
  Stream2Mmap_12__ap_done,
  Stream2Mmap_12__ap_idle,
  Stream2Mmap_13___n__q0,
  Stream2Mmap_13___rmem13__q0,
  Stream2Mmap_13__ap_start,
  Stream2Mmap_13__ap_ready,
  Stream2Mmap_13__ap_done,
  Stream2Mmap_13__ap_idle,
  Stream2Mmap_14___n__q0,
  Stream2Mmap_14___rmem14__q0,
  Stream2Mmap_14__ap_start,
  Stream2Mmap_14__ap_ready,
  Stream2Mmap_14__ap_done,
  Stream2Mmap_14__ap_idle,
  Stream2Mmap_15___n__q0,
  Stream2Mmap_15___rmem15__q0,
  Stream2Mmap_15__ap_start,
  Stream2Mmap_15__ap_ready,
  Stream2Mmap_15__ap_done,
  Stream2Mmap_15__ap_idle,
  Stream2Mmap_16___n__q0,
  Stream2Mmap_16___rmem16__q0,
  Stream2Mmap_16__ap_start,
  Stream2Mmap_16__ap_ready,
  Stream2Mmap_16__ap_done,
  Stream2Mmap_16__ap_idle,
  Stream2Mmap_17___n__q0,
  Stream2Mmap_17___rmem17__q0,
  Stream2Mmap_17__ap_start,
  Stream2Mmap_17__ap_ready,
  Stream2Mmap_17__ap_done,
  Stream2Mmap_17__ap_idle,
  Stream2Mmap_18___n__q0,
  Stream2Mmap_18___rmem18__q0,
  Stream2Mmap_18__ap_start,
  Stream2Mmap_18__ap_ready,
  Stream2Mmap_18__ap_done,
  Stream2Mmap_18__ap_idle,
  Stream2Mmap_19___n__q0,
  Stream2Mmap_19___rmem19__q0,
  Stream2Mmap_19__ap_start,
  Stream2Mmap_19__ap_ready,
  Stream2Mmap_19__ap_done,
  Stream2Mmap_19__ap_idle,
  Stream2Mmap_20___n__q0,
  Stream2Mmap_20___rmem20__q0,
  Stream2Mmap_20__ap_start,
  Stream2Mmap_20__ap_ready,
  Stream2Mmap_20__ap_done,
  Stream2Mmap_20__ap_idle,
  Stream2Mmap_21___n__q0,
  Stream2Mmap_21___rmem21__q0,
  Stream2Mmap_21__ap_start,
  Stream2Mmap_21__ap_ready,
  Stream2Mmap_21__ap_done,
  Stream2Mmap_21__ap_idle,
  Stream2Mmap_22___n__q0,
  Stream2Mmap_22___rmem22__q0,
  Stream2Mmap_22__ap_start,
  Stream2Mmap_22__ap_ready,
  Stream2Mmap_22__ap_done,
  Stream2Mmap_22__ap_idle,
  Stream2Mmap_23___n__q0,
  Stream2Mmap_23___rmem23__q0,
  Stream2Mmap_23__ap_start,
  Stream2Mmap_23__ap_ready,
  Stream2Mmap_23__ap_done,
  Stream2Mmap_23__ap_idle,
  Stream2Mmap_24___n__q0,
  Stream2Mmap_24___rmem24__q0,
  Stream2Mmap_24__ap_start,
  Stream2Mmap_24__ap_ready,
  Stream2Mmap_24__ap_done,
  Stream2Mmap_24__ap_idle,
  Stream2Mmap_25___n__q0,
  Stream2Mmap_25___rmem25__q0,
  Stream2Mmap_25__ap_start,
  Stream2Mmap_25__ap_ready,
  Stream2Mmap_25__ap_done,
  Stream2Mmap_25__ap_idle,
  Stream2Mmap_26___n__q0,
  Stream2Mmap_26___rmem26__q0,
  Stream2Mmap_26__ap_start,
  Stream2Mmap_26__ap_ready,
  Stream2Mmap_26__ap_done,
  Stream2Mmap_26__ap_idle,
  yshift_0___n__q0,
  yshift_0__ap_start,
  yshift_0__ap_ready,
  yshift_0__ap_done,
  yshift_0__ap_idle,
  yshift_1___n__q0,
  yshift_1__ap_start,
  yshift_1__ap_ready,
  yshift_1__ap_done,
  yshift_1__ap_idle,
  yshift_2___n__q0,
  yshift_2__ap_start,
  yshift_2__ap_ready,
  yshift_2__ap_done,
  yshift_2__ap_idle,
  yshift_3___n__q0,
  yshift_3__ap_start,
  yshift_3__ap_ready,
  yshift_3__ap_done,
  yshift_3__ap_idle,
  yshift_4___n__q0,
  yshift_4__ap_start,
  yshift_4__ap_ready,
  yshift_4__ap_done,
  yshift_4__ap_idle,
  yshift_5___n__q0,
  yshift_5__ap_start,
  yshift_5__ap_ready,
  yshift_5__ap_done,
  yshift_5__ap_idle,
  yshift_6___n__q0,
  yshift_6__ap_start,
  yshift_6__ap_ready,
  yshift_6__ap_done,
  yshift_6__ap_idle,
  yshift_7___n__q0,
  yshift_7__ap_start,
  yshift_7__ap_ready,
  yshift_7__ap_done,
  yshift_7__ap_idle,
  yshift_8___n__q0,
  yshift_8__ap_start,
  yshift_8__ap_ready,
  yshift_8__ap_done,
  yshift_8__ap_idle,
  yshift_9___n__q0,
  yshift_9__ap_start,
  yshift_9__ap_ready,
  yshift_9__ap_done,
  yshift_9__ap_idle,
  yshift_10___n__q0,
  yshift_10__ap_start,
  yshift_10__ap_ready,
  yshift_10__ap_done,
  yshift_10__ap_idle,
  yshift_11___n__q0,
  yshift_11__ap_start,
  yshift_11__ap_ready,
  yshift_11__ap_done,
  yshift_11__ap_idle,
  yshift_12___n__q0,
  yshift_12__ap_start,
  yshift_12__ap_ready,
  yshift_12__ap_done,
  yshift_12__ap_idle,
  yshift_13___n__q0,
  yshift_13__ap_start,
  yshift_13__ap_ready,
  yshift_13__ap_done,
  yshift_13__ap_idle,
  yshift_14___n__q0,
  yshift_14__ap_start,
  yshift_14__ap_ready,
  yshift_14__ap_done,
  yshift_14__ap_idle,
  yshift_15___n__q0,
  yshift_15__ap_start,
  yshift_15__ap_ready,
  yshift_15__ap_done,
  yshift_15__ap_idle,
  yshift_16___n__q0,
  yshift_16__ap_start,
  yshift_16__ap_ready,
  yshift_16__ap_done,
  yshift_16__ap_idle,
  yshift_17___n__q0,
  yshift_17__ap_start,
  yshift_17__ap_ready,
  yshift_17__ap_done,
  yshift_17__ap_idle,
  yshift_18___n__q0,
  yshift_18__ap_start,
  yshift_18__ap_ready,
  yshift_18__ap_done,
  yshift_18__ap_idle,
  yshift_19___n__q0,
  yshift_19__ap_start,
  yshift_19__ap_ready,
  yshift_19__ap_done,
  yshift_19__ap_idle,
  yshift_20___n__q0,
  yshift_20__ap_start,
  yshift_20__ap_ready,
  yshift_20__ap_done,
  yshift_20__ap_idle,
  yshift_21___n__q0,
  yshift_21__ap_start,
  yshift_21__ap_ready,
  yshift_21__ap_done,
  yshift_21__ap_idle,
  yshift_22___n__q0,
  yshift_22__ap_start,
  yshift_22__ap_ready,
  yshift_22__ap_done,
  yshift_22__ap_idle,
  yshift_23___n__q0,
  yshift_23__ap_start,
  yshift_23__ap_ready,
  yshift_23__ap_done,
  yshift_23__ap_idle,
  yshift_24___n__q0,
  yshift_24__ap_start,
  yshift_24__ap_ready,
  yshift_24__ap_done,
  yshift_24__ap_idle,
  yshift_25___n__q0,
  yshift_25__ap_start,
  yshift_25__ap_ready,
  yshift_25__ap_done,
  yshift_25__ap_idle,
  yshift_26___n__q0,
  yshift_26__ap_start,
  yshift_26__ap_ready,
  yshift_26__ap_done,
  yshift_26__ap_idle
);

  // pragma RS clk port=ap_clk
  // pragma RS rst port=ap_rst_n active=low
  // pragma RS ap-ctrl ap_start=ap_start ap_done=ap_done ap_idle=ap_idle ap_ready=ap_ready scalar=(rmem0|rmem1|rmem2|rmem3|rmem4|rmem5|rmem6|rmem7|rmem8|rmem9|rmem10|rmem11|rmem12|rmem13|rmem14|rmem15|rmem16|rmem17|rmem18|rmem19|rmem20|rmem21|rmem22|rmem23|rmem24|rmem25|rmem26|n)
  // pragma RS ap-ctrl ap_start=Mmap2Stream_0__ap_start ap_done=Mmap2Stream_0__ap_done ap_idle=Mmap2Stream_0__ap_idle ap_ready=Mmap2Stream_0__ap_ready scalar=Mmap2Stream_0___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_1__ap_start ap_done=Mmap2Stream_1__ap_done ap_idle=Mmap2Stream_1__ap_idle ap_ready=Mmap2Stream_1__ap_ready scalar=Mmap2Stream_1___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_2__ap_start ap_done=Mmap2Stream_2__ap_done ap_idle=Mmap2Stream_2__ap_idle ap_ready=Mmap2Stream_2__ap_ready scalar=Mmap2Stream_2___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_3__ap_start ap_done=Mmap2Stream_3__ap_done ap_idle=Mmap2Stream_3__ap_idle ap_ready=Mmap2Stream_3__ap_ready scalar=Mmap2Stream_3___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_4__ap_start ap_done=Mmap2Stream_4__ap_done ap_idle=Mmap2Stream_4__ap_idle ap_ready=Mmap2Stream_4__ap_ready scalar=Mmap2Stream_4___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_5__ap_start ap_done=Mmap2Stream_5__ap_done ap_idle=Mmap2Stream_5__ap_idle ap_ready=Mmap2Stream_5__ap_ready scalar=Mmap2Stream_5___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_6__ap_start ap_done=Mmap2Stream_6__ap_done ap_idle=Mmap2Stream_6__ap_idle ap_ready=Mmap2Stream_6__ap_ready scalar=Mmap2Stream_6___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_7__ap_start ap_done=Mmap2Stream_7__ap_done ap_idle=Mmap2Stream_7__ap_idle ap_ready=Mmap2Stream_7__ap_ready scalar=Mmap2Stream_7___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_8__ap_start ap_done=Mmap2Stream_8__ap_done ap_idle=Mmap2Stream_8__ap_idle ap_ready=Mmap2Stream_8__ap_ready scalar=Mmap2Stream_8___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_9__ap_start ap_done=Mmap2Stream_9__ap_done ap_idle=Mmap2Stream_9__ap_idle ap_ready=Mmap2Stream_9__ap_ready scalar=Mmap2Stream_9___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_10__ap_start ap_done=Mmap2Stream_10__ap_done ap_idle=Mmap2Stream_10__ap_idle ap_ready=Mmap2Stream_10__ap_ready scalar=Mmap2Stream_10___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_11__ap_start ap_done=Mmap2Stream_11__ap_done ap_idle=Mmap2Stream_11__ap_idle ap_ready=Mmap2Stream_11__ap_ready scalar=Mmap2Stream_11___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_12__ap_start ap_done=Mmap2Stream_12__ap_done ap_idle=Mmap2Stream_12__ap_idle ap_ready=Mmap2Stream_12__ap_ready scalar=Mmap2Stream_12___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_13__ap_start ap_done=Mmap2Stream_13__ap_done ap_idle=Mmap2Stream_13__ap_idle ap_ready=Mmap2Stream_13__ap_ready scalar=Mmap2Stream_13___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_14__ap_start ap_done=Mmap2Stream_14__ap_done ap_idle=Mmap2Stream_14__ap_idle ap_ready=Mmap2Stream_14__ap_ready scalar=Mmap2Stream_14___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_15__ap_start ap_done=Mmap2Stream_15__ap_done ap_idle=Mmap2Stream_15__ap_idle ap_ready=Mmap2Stream_15__ap_ready scalar=Mmap2Stream_15___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_16__ap_start ap_done=Mmap2Stream_16__ap_done ap_idle=Mmap2Stream_16__ap_idle ap_ready=Mmap2Stream_16__ap_ready scalar=Mmap2Stream_16___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_17__ap_start ap_done=Mmap2Stream_17__ap_done ap_idle=Mmap2Stream_17__ap_idle ap_ready=Mmap2Stream_17__ap_ready scalar=Mmap2Stream_17___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_18__ap_start ap_done=Mmap2Stream_18__ap_done ap_idle=Mmap2Stream_18__ap_idle ap_ready=Mmap2Stream_18__ap_ready scalar=Mmap2Stream_18___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_19__ap_start ap_done=Mmap2Stream_19__ap_done ap_idle=Mmap2Stream_19__ap_idle ap_ready=Mmap2Stream_19__ap_ready scalar=Mmap2Stream_19___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_20__ap_start ap_done=Mmap2Stream_20__ap_done ap_idle=Mmap2Stream_20__ap_idle ap_ready=Mmap2Stream_20__ap_ready scalar=Mmap2Stream_20___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_21__ap_start ap_done=Mmap2Stream_21__ap_done ap_idle=Mmap2Stream_21__ap_idle ap_ready=Mmap2Stream_21__ap_ready scalar=Mmap2Stream_21___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_22__ap_start ap_done=Mmap2Stream_22__ap_done ap_idle=Mmap2Stream_22__ap_idle ap_ready=Mmap2Stream_22__ap_ready scalar=Mmap2Stream_22___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_23__ap_start ap_done=Mmap2Stream_23__ap_done ap_idle=Mmap2Stream_23__ap_idle ap_ready=Mmap2Stream_23__ap_ready scalar=Mmap2Stream_23___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_24__ap_start ap_done=Mmap2Stream_24__ap_done ap_idle=Mmap2Stream_24__ap_idle ap_ready=Mmap2Stream_24__ap_ready scalar=Mmap2Stream_24___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_25__ap_start ap_done=Mmap2Stream_25__ap_done ap_idle=Mmap2Stream_25__ap_idle ap_ready=Mmap2Stream_25__ap_ready scalar=Mmap2Stream_25___.*
  // pragma RS ap-ctrl ap_start=Mmap2Stream_26__ap_start ap_done=Mmap2Stream_26__ap_done ap_idle=Mmap2Stream_26__ap_idle ap_ready=Mmap2Stream_26__ap_ready scalar=Mmap2Stream_26___.*
  // pragma RS ap-ctrl ap_start=Stream2Mmap_0__ap_start ap_done=Stream2Mmap_0__ap_done ap_idle=Stream2Mmap_0__ap_idle ap_ready=Stream2Mmap_0__ap_ready scalar=Stream2Mmap_0___.*
  // pragma RS ap-ctrl ap_start=Stream2Mmap_1__ap_start ap_done=Stream2Mmap_1__ap_done ap_idle=Stream2Mmap_1__ap_idle ap_ready=Stream2Mmap_1__ap_ready scalar=Stream2Mmap_1___.*
  // pragma RS ap-ctrl ap_start=Stream2Mmap_2__ap_start ap_done=Stream2Mmap_2__ap_done ap_idle=Stream2Mmap_2__ap_idle ap_ready=Stream2Mmap_2__ap_ready scalar=Stream2Mmap_2___.*
  // pragma RS ap-ctrl ap_start=Stream2Mmap_3__ap_start ap_done=Stream2Mmap_3__ap_done ap_idle=Stream2Mmap_3__ap_idle ap_ready=Stream2Mmap_3__ap_ready scalar=Stream2Mmap_3___.*
  // pragma RS ap-ctrl ap_start=Stream2Mmap_4__ap_start ap_done=Stream2Mmap_4__ap_done ap_idle=Stream2Mmap_4__ap_idle ap_ready=Stream2Mmap_4__ap_ready scalar=Stream2Mmap_4___.*
  // pragma RS ap-ctrl ap_start=Stream2Mmap_5__ap_start ap_done=Stream2Mmap_5__ap_done ap_idle=Stream2Mmap_5__ap_idle ap_ready=Stream2Mmap_5__ap_ready scalar=Stream2Mmap_5___.*
  // pragma RS ap-ctrl ap_start=Stream2Mmap_6__ap_start ap_done=Stream2Mmap_6__ap_done ap_idle=Stream2Mmap_6__ap_idle ap_ready=Stream2Mmap_6__ap_ready scalar=Stream2Mmap_6___.*
  // pragma RS ap-ctrl ap_start=Stream2Mmap_7__ap_start ap_done=Stream2Mmap_7__ap_done ap_idle=Stream2Mmap_7__ap_idle ap_ready=Stream2Mmap_7__ap_ready scalar=Stream2Mmap_7___.*
  // pragma RS ap-ctrl ap_start=Stream2Mmap_8__ap_start ap_done=Stream2Mmap_8__ap_done ap_idle=Stream2Mmap_8__ap_idle ap_ready=Stream2Mmap_8__ap_ready scalar=Stream2Mmap_8___.*
  // pragma RS ap-ctrl ap_start=Stream2Mmap_9__ap_start ap_done=Stream2Mmap_9__ap_done ap_idle=Stream2Mmap_9__ap_idle ap_ready=Stream2Mmap_9__ap_ready scalar=Stream2Mmap_9___.*
  // pragma RS ap-ctrl ap_start=Stream2Mmap_10__ap_start ap_done=Stream2Mmap_10__ap_done ap_idle=Stream2Mmap_10__ap_idle ap_ready=Stream2Mmap_10__ap_ready scalar=Stream2Mmap_10___.*
  // pragma RS ap-ctrl ap_start=Stream2Mmap_11__ap_start ap_done=Stream2Mmap_11__ap_done ap_idle=Stream2Mmap_11__ap_idle ap_ready=Stream2Mmap_11__ap_ready scalar=Stream2Mmap_11___.*
  // pragma RS ap-ctrl ap_start=Stream2Mmap_12__ap_start ap_done=Stream2Mmap_12__ap_done ap_idle=Stream2Mmap_12__ap_idle ap_ready=Stream2Mmap_12__ap_ready scalar=Stream2Mmap_12___.*
  // pragma RS ap-ctrl ap_start=Stream2Mmap_13__ap_start ap_done=Stream2Mmap_13__ap_done ap_idle=Stream2Mmap_13__ap_idle ap_ready=Stream2Mmap_13__ap_ready scalar=Stream2Mmap_13___.*
  // pragma RS ap-ctrl ap_start=Stream2Mmap_14__ap_start ap_done=Stream2Mmap_14__ap_done ap_idle=Stream2Mmap_14__ap_idle ap_ready=Stream2Mmap_14__ap_ready scalar=Stream2Mmap_14___.*
  // pragma RS ap-ctrl ap_start=Stream2Mmap_15__ap_start ap_done=Stream2Mmap_15__ap_done ap_idle=Stream2Mmap_15__ap_idle ap_ready=Stream2Mmap_15__ap_ready scalar=Stream2Mmap_15___.*
  // pragma RS ap-ctrl ap_start=Stream2Mmap_16__ap_start ap_done=Stream2Mmap_16__ap_done ap_idle=Stream2Mmap_16__ap_idle ap_ready=Stream2Mmap_16__ap_ready scalar=Stream2Mmap_16___.*
  // pragma RS ap-ctrl ap_start=Stream2Mmap_17__ap_start ap_done=Stream2Mmap_17__ap_done ap_idle=Stream2Mmap_17__ap_idle ap_ready=Stream2Mmap_17__ap_ready scalar=Stream2Mmap_17___.*
  // pragma RS ap-ctrl ap_start=Stream2Mmap_18__ap_start ap_done=Stream2Mmap_18__ap_done ap_idle=Stream2Mmap_18__ap_idle ap_ready=Stream2Mmap_18__ap_ready scalar=Stream2Mmap_18___.*
  // pragma RS ap-ctrl ap_start=Stream2Mmap_19__ap_start ap_done=Stream2Mmap_19__ap_done ap_idle=Stream2Mmap_19__ap_idle ap_ready=Stream2Mmap_19__ap_ready scalar=Stream2Mmap_19___.*
  // pragma RS ap-ctrl ap_start=Stream2Mmap_20__ap_start ap_done=Stream2Mmap_20__ap_done ap_idle=Stream2Mmap_20__ap_idle ap_ready=Stream2Mmap_20__ap_ready scalar=Stream2Mmap_20___.*
  // pragma RS ap-ctrl ap_start=Stream2Mmap_21__ap_start ap_done=Stream2Mmap_21__ap_done ap_idle=Stream2Mmap_21__ap_idle ap_ready=Stream2Mmap_21__ap_ready scalar=Stream2Mmap_21___.*
  // pragma RS ap-ctrl ap_start=Stream2Mmap_22__ap_start ap_done=Stream2Mmap_22__ap_done ap_idle=Stream2Mmap_22__ap_idle ap_ready=Stream2Mmap_22__ap_ready scalar=Stream2Mmap_22___.*
  // pragma RS ap-ctrl ap_start=Stream2Mmap_23__ap_start ap_done=Stream2Mmap_23__ap_done ap_idle=Stream2Mmap_23__ap_idle ap_ready=Stream2Mmap_23__ap_ready scalar=Stream2Mmap_23___.*
  // pragma RS ap-ctrl ap_start=Stream2Mmap_24__ap_start ap_done=Stream2Mmap_24__ap_done ap_idle=Stream2Mmap_24__ap_idle ap_ready=Stream2Mmap_24__ap_ready scalar=Stream2Mmap_24___.*
  // pragma RS ap-ctrl ap_start=Stream2Mmap_25__ap_start ap_done=Stream2Mmap_25__ap_done ap_idle=Stream2Mmap_25__ap_idle ap_ready=Stream2Mmap_25__ap_ready scalar=Stream2Mmap_25___.*
  // pragma RS ap-ctrl ap_start=Stream2Mmap_26__ap_start ap_done=Stream2Mmap_26__ap_done ap_idle=Stream2Mmap_26__ap_idle ap_ready=Stream2Mmap_26__ap_ready scalar=Stream2Mmap_26___.*
  // pragma RS ap-ctrl ap_start=yshift_0__ap_start ap_done=yshift_0__ap_done ap_idle=yshift_0__ap_idle ap_ready=yshift_0__ap_ready scalar=yshift_0___.*
  // pragma RS ap-ctrl ap_start=yshift_1__ap_start ap_done=yshift_1__ap_done ap_idle=yshift_1__ap_idle ap_ready=yshift_1__ap_ready scalar=yshift_1___.*
  // pragma RS ap-ctrl ap_start=yshift_2__ap_start ap_done=yshift_2__ap_done ap_idle=yshift_2__ap_idle ap_ready=yshift_2__ap_ready scalar=yshift_2___.*
  // pragma RS ap-ctrl ap_start=yshift_3__ap_start ap_done=yshift_3__ap_done ap_idle=yshift_3__ap_idle ap_ready=yshift_3__ap_ready scalar=yshift_3___.*
  // pragma RS ap-ctrl ap_start=yshift_4__ap_start ap_done=yshift_4__ap_done ap_idle=yshift_4__ap_idle ap_ready=yshift_4__ap_ready scalar=yshift_4___.*
  // pragma RS ap-ctrl ap_start=yshift_5__ap_start ap_done=yshift_5__ap_done ap_idle=yshift_5__ap_idle ap_ready=yshift_5__ap_ready scalar=yshift_5___.*
  // pragma RS ap-ctrl ap_start=yshift_6__ap_start ap_done=yshift_6__ap_done ap_idle=yshift_6__ap_idle ap_ready=yshift_6__ap_ready scalar=yshift_6___.*
  // pragma RS ap-ctrl ap_start=yshift_7__ap_start ap_done=yshift_7__ap_done ap_idle=yshift_7__ap_idle ap_ready=yshift_7__ap_ready scalar=yshift_7___.*
  // pragma RS ap-ctrl ap_start=yshift_8__ap_start ap_done=yshift_8__ap_done ap_idle=yshift_8__ap_idle ap_ready=yshift_8__ap_ready scalar=yshift_8___.*
  // pragma RS ap-ctrl ap_start=yshift_9__ap_start ap_done=yshift_9__ap_done ap_idle=yshift_9__ap_idle ap_ready=yshift_9__ap_ready scalar=yshift_9___.*
  // pragma RS ap-ctrl ap_start=yshift_10__ap_start ap_done=yshift_10__ap_done ap_idle=yshift_10__ap_idle ap_ready=yshift_10__ap_ready scalar=yshift_10___.*
  // pragma RS ap-ctrl ap_start=yshift_11__ap_start ap_done=yshift_11__ap_done ap_idle=yshift_11__ap_idle ap_ready=yshift_11__ap_ready scalar=yshift_11___.*
  // pragma RS ap-ctrl ap_start=yshift_12__ap_start ap_done=yshift_12__ap_done ap_idle=yshift_12__ap_idle ap_ready=yshift_12__ap_ready scalar=yshift_12___.*
  // pragma RS ap-ctrl ap_start=yshift_13__ap_start ap_done=yshift_13__ap_done ap_idle=yshift_13__ap_idle ap_ready=yshift_13__ap_ready scalar=yshift_13___.*
  // pragma RS ap-ctrl ap_start=yshift_14__ap_start ap_done=yshift_14__ap_done ap_idle=yshift_14__ap_idle ap_ready=yshift_14__ap_ready scalar=yshift_14___.*
  // pragma RS ap-ctrl ap_start=yshift_15__ap_start ap_done=yshift_15__ap_done ap_idle=yshift_15__ap_idle ap_ready=yshift_15__ap_ready scalar=yshift_15___.*
  // pragma RS ap-ctrl ap_start=yshift_16__ap_start ap_done=yshift_16__ap_done ap_idle=yshift_16__ap_idle ap_ready=yshift_16__ap_ready scalar=yshift_16___.*
  // pragma RS ap-ctrl ap_start=yshift_17__ap_start ap_done=yshift_17__ap_done ap_idle=yshift_17__ap_idle ap_ready=yshift_17__ap_ready scalar=yshift_17___.*
  // pragma RS ap-ctrl ap_start=yshift_18__ap_start ap_done=yshift_18__ap_done ap_idle=yshift_18__ap_idle ap_ready=yshift_18__ap_ready scalar=yshift_18___.*
  // pragma RS ap-ctrl ap_start=yshift_19__ap_start ap_done=yshift_19__ap_done ap_idle=yshift_19__ap_idle ap_ready=yshift_19__ap_ready scalar=yshift_19___.*
  // pragma RS ap-ctrl ap_start=yshift_20__ap_start ap_done=yshift_20__ap_done ap_idle=yshift_20__ap_idle ap_ready=yshift_20__ap_ready scalar=yshift_20___.*
  // pragma RS ap-ctrl ap_start=yshift_21__ap_start ap_done=yshift_21__ap_done ap_idle=yshift_21__ap_idle ap_ready=yshift_21__ap_ready scalar=yshift_21___.*
  // pragma RS ap-ctrl ap_start=yshift_22__ap_start ap_done=yshift_22__ap_done ap_idle=yshift_22__ap_idle ap_ready=yshift_22__ap_ready scalar=yshift_22___.*
  // pragma RS ap-ctrl ap_start=yshift_23__ap_start ap_done=yshift_23__ap_done ap_idle=yshift_23__ap_idle ap_ready=yshift_23__ap_ready scalar=yshift_23___.*
  // pragma RS ap-ctrl ap_start=yshift_24__ap_start ap_done=yshift_24__ap_done ap_idle=yshift_24__ap_idle ap_ready=yshift_24__ap_ready scalar=yshift_24___.*
  // pragma RS ap-ctrl ap_start=yshift_25__ap_start ap_done=yshift_25__ap_done ap_idle=yshift_25__ap_idle ap_ready=yshift_25__ap_ready scalar=yshift_25___.*
  // pragma RS ap-ctrl ap_start=yshift_26__ap_start ap_done=yshift_26__ap_done ap_idle=yshift_26__ap_idle ap_ready=yshift_26__ap_ready scalar=yshift_26___.*

  input ap_clk;
  input ap_rst_n;
  input ap_start;
  output ap_ready;
  output ap_done;
  output ap_idle;
  input [63:0] n;
  input [63:0] rmem0;
  input [63:0] rmem1;
  input [63:0] rmem2;
  input [63:0] rmem3;
  input [63:0] rmem4;
  input [63:0] rmem5;
  input [63:0] rmem6;
  input [63:0] rmem7;
  input [63:0] rmem8;
  input [63:0] rmem9;
  input [63:0] rmem10;
  input [63:0] rmem11;
  input [63:0] rmem12;
  input [63:0] rmem13;
  input [63:0] rmem14;
  input [63:0] rmem15;
  input [63:0] rmem16;
  input [63:0] rmem17;
  input [63:0] rmem18;
  input [63:0] rmem19;
  input [63:0] rmem20;
  input [63:0] rmem21;
  input [63:0] rmem22;
  input [63:0] rmem23;
  input [63:0] rmem24;
  input [63:0] rmem25;
  input [63:0] rmem26;
  output [63:0] Mmap2Stream_0___n__q0;
  output [63:0] Mmap2Stream_0___rmem0__q0;
  output Mmap2Stream_0__ap_start;
  input Mmap2Stream_0__ap_ready;
  input Mmap2Stream_0__ap_done;
  input Mmap2Stream_0__ap_idle;
  output [63:0] Mmap2Stream_1___n__q0;
  output [63:0] Mmap2Stream_1___rmem1__q0;
  output Mmap2Stream_1__ap_start;
  input Mmap2Stream_1__ap_ready;
  input Mmap2Stream_1__ap_done;
  input Mmap2Stream_1__ap_idle;
  output [63:0] Mmap2Stream_2___n__q0;
  output [63:0] Mmap2Stream_2___rmem2__q0;
  output Mmap2Stream_2__ap_start;
  input Mmap2Stream_2__ap_ready;
  input Mmap2Stream_2__ap_done;
  input Mmap2Stream_2__ap_idle;
  output [63:0] Mmap2Stream_3___n__q0;
  output [63:0] Mmap2Stream_3___rmem3__q0;
  output Mmap2Stream_3__ap_start;
  input Mmap2Stream_3__ap_ready;
  input Mmap2Stream_3__ap_done;
  input Mmap2Stream_3__ap_idle;
  output [63:0] Mmap2Stream_4___n__q0;
  output [63:0] Mmap2Stream_4___rmem4__q0;
  output Mmap2Stream_4__ap_start;
  input Mmap2Stream_4__ap_ready;
  input Mmap2Stream_4__ap_done;
  input Mmap2Stream_4__ap_idle;
  output [63:0] Mmap2Stream_5___n__q0;
  output [63:0] Mmap2Stream_5___rmem5__q0;
  output Mmap2Stream_5__ap_start;
  input Mmap2Stream_5__ap_ready;
  input Mmap2Stream_5__ap_done;
  input Mmap2Stream_5__ap_idle;
  output [63:0] Mmap2Stream_6___n__q0;
  output [63:0] Mmap2Stream_6___rmem6__q0;
  output Mmap2Stream_6__ap_start;
  input Mmap2Stream_6__ap_ready;
  input Mmap2Stream_6__ap_done;
  input Mmap2Stream_6__ap_idle;
  output [63:0] Mmap2Stream_7___n__q0;
  output [63:0] Mmap2Stream_7___rmem7__q0;
  output Mmap2Stream_7__ap_start;
  input Mmap2Stream_7__ap_ready;
  input Mmap2Stream_7__ap_done;
  input Mmap2Stream_7__ap_idle;
  output [63:0] Mmap2Stream_8___n__q0;
  output [63:0] Mmap2Stream_8___rmem8__q0;
  output Mmap2Stream_8__ap_start;
  input Mmap2Stream_8__ap_ready;
  input Mmap2Stream_8__ap_done;
  input Mmap2Stream_8__ap_idle;
  output [63:0] Mmap2Stream_9___n__q0;
  output [63:0] Mmap2Stream_9___rmem9__q0;
  output Mmap2Stream_9__ap_start;
  input Mmap2Stream_9__ap_ready;
  input Mmap2Stream_9__ap_done;
  input Mmap2Stream_9__ap_idle;
  output [63:0] Mmap2Stream_10___n__q0;
  output [63:0] Mmap2Stream_10___rmem10__q0;
  output Mmap2Stream_10__ap_start;
  input Mmap2Stream_10__ap_ready;
  input Mmap2Stream_10__ap_done;
  input Mmap2Stream_10__ap_idle;
  output [63:0] Mmap2Stream_11___n__q0;
  output [63:0] Mmap2Stream_11___rmem11__q0;
  output Mmap2Stream_11__ap_start;
  input Mmap2Stream_11__ap_ready;
  input Mmap2Stream_11__ap_done;
  input Mmap2Stream_11__ap_idle;
  output [63:0] Mmap2Stream_12___n__q0;
  output [63:0] Mmap2Stream_12___rmem12__q0;
  output Mmap2Stream_12__ap_start;
  input Mmap2Stream_12__ap_ready;
  input Mmap2Stream_12__ap_done;
  input Mmap2Stream_12__ap_idle;
  output [63:0] Mmap2Stream_13___n__q0;
  output [63:0] Mmap2Stream_13___rmem13__q0;
  output Mmap2Stream_13__ap_start;
  input Mmap2Stream_13__ap_ready;
  input Mmap2Stream_13__ap_done;
  input Mmap2Stream_13__ap_idle;
  output [63:0] Mmap2Stream_14___n__q0;
  output [63:0] Mmap2Stream_14___rmem14__q0;
  output Mmap2Stream_14__ap_start;
  input Mmap2Stream_14__ap_ready;
  input Mmap2Stream_14__ap_done;
  input Mmap2Stream_14__ap_idle;
  output [63:0] Mmap2Stream_15___n__q0;
  output [63:0] Mmap2Stream_15___rmem15__q0;
  output Mmap2Stream_15__ap_start;
  input Mmap2Stream_15__ap_ready;
  input Mmap2Stream_15__ap_done;
  input Mmap2Stream_15__ap_idle;
  output [63:0] Mmap2Stream_16___n__q0;
  output [63:0] Mmap2Stream_16___rmem16__q0;
  output Mmap2Stream_16__ap_start;
  input Mmap2Stream_16__ap_ready;
  input Mmap2Stream_16__ap_done;
  input Mmap2Stream_16__ap_idle;
  output [63:0] Mmap2Stream_17___n__q0;
  output [63:0] Mmap2Stream_17___rmem17__q0;
  output Mmap2Stream_17__ap_start;
  input Mmap2Stream_17__ap_ready;
  input Mmap2Stream_17__ap_done;
  input Mmap2Stream_17__ap_idle;
  output [63:0] Mmap2Stream_18___n__q0;
  output [63:0] Mmap2Stream_18___rmem18__q0;
  output Mmap2Stream_18__ap_start;
  input Mmap2Stream_18__ap_ready;
  input Mmap2Stream_18__ap_done;
  input Mmap2Stream_18__ap_idle;
  output [63:0] Mmap2Stream_19___n__q0;
  output [63:0] Mmap2Stream_19___rmem19__q0;
  output Mmap2Stream_19__ap_start;
  input Mmap2Stream_19__ap_ready;
  input Mmap2Stream_19__ap_done;
  input Mmap2Stream_19__ap_idle;
  output [63:0] Mmap2Stream_20___n__q0;
  output [63:0] Mmap2Stream_20___rmem20__q0;
  output Mmap2Stream_20__ap_start;
  input Mmap2Stream_20__ap_ready;
  input Mmap2Stream_20__ap_done;
  input Mmap2Stream_20__ap_idle;
  output [63:0] Mmap2Stream_21___n__q0;
  output [63:0] Mmap2Stream_21___rmem21__q0;
  output Mmap2Stream_21__ap_start;
  input Mmap2Stream_21__ap_ready;
  input Mmap2Stream_21__ap_done;
  input Mmap2Stream_21__ap_idle;
  output [63:0] Mmap2Stream_22___n__q0;
  output [63:0] Mmap2Stream_22___rmem22__q0;
  output Mmap2Stream_22__ap_start;
  input Mmap2Stream_22__ap_ready;
  input Mmap2Stream_22__ap_done;
  input Mmap2Stream_22__ap_idle;
  output [63:0] Mmap2Stream_23___n__q0;
  output [63:0] Mmap2Stream_23___rmem23__q0;
  output Mmap2Stream_23__ap_start;
  input Mmap2Stream_23__ap_ready;
  input Mmap2Stream_23__ap_done;
  input Mmap2Stream_23__ap_idle;
  output [63:0] Mmap2Stream_24___n__q0;
  output [63:0] Mmap2Stream_24___rmem24__q0;
  output Mmap2Stream_24__ap_start;
  input Mmap2Stream_24__ap_ready;
  input Mmap2Stream_24__ap_done;
  input Mmap2Stream_24__ap_idle;
  output [63:0] Mmap2Stream_25___n__q0;
  output [63:0] Mmap2Stream_25___rmem25__q0;
  output Mmap2Stream_25__ap_start;
  input Mmap2Stream_25__ap_ready;
  input Mmap2Stream_25__ap_done;
  input Mmap2Stream_25__ap_idle;
  output [63:0] Mmap2Stream_26___n__q0;
  output [63:0] Mmap2Stream_26___rmem26__q0;
  output Mmap2Stream_26__ap_start;
  input Mmap2Stream_26__ap_ready;
  input Mmap2Stream_26__ap_done;
  input Mmap2Stream_26__ap_idle;
  output [63:0] Stream2Mmap_0___n__q0;
  output [63:0] Stream2Mmap_0___rmem0__q0;
  output Stream2Mmap_0__ap_start;
  input Stream2Mmap_0__ap_ready;
  input Stream2Mmap_0__ap_done;
  input Stream2Mmap_0__ap_idle;
  output [63:0] Stream2Mmap_1___n__q0;
  output [63:0] Stream2Mmap_1___rmem1__q0;
  output Stream2Mmap_1__ap_start;
  input Stream2Mmap_1__ap_ready;
  input Stream2Mmap_1__ap_done;
  input Stream2Mmap_1__ap_idle;
  output [63:0] Stream2Mmap_2___n__q0;
  output [63:0] Stream2Mmap_2___rmem2__q0;
  output Stream2Mmap_2__ap_start;
  input Stream2Mmap_2__ap_ready;
  input Stream2Mmap_2__ap_done;
  input Stream2Mmap_2__ap_idle;
  output [63:0] Stream2Mmap_3___n__q0;
  output [63:0] Stream2Mmap_3___rmem3__q0;
  output Stream2Mmap_3__ap_start;
  input Stream2Mmap_3__ap_ready;
  input Stream2Mmap_3__ap_done;
  input Stream2Mmap_3__ap_idle;
  output [63:0] Stream2Mmap_4___n__q0;
  output [63:0] Stream2Mmap_4___rmem4__q0;
  output Stream2Mmap_4__ap_start;
  input Stream2Mmap_4__ap_ready;
  input Stream2Mmap_4__ap_done;
  input Stream2Mmap_4__ap_idle;
  output [63:0] Stream2Mmap_5___n__q0;
  output [63:0] Stream2Mmap_5___rmem5__q0;
  output Stream2Mmap_5__ap_start;
  input Stream2Mmap_5__ap_ready;
  input Stream2Mmap_5__ap_done;
  input Stream2Mmap_5__ap_idle;
  output [63:0] Stream2Mmap_6___n__q0;
  output [63:0] Stream2Mmap_6___rmem6__q0;
  output Stream2Mmap_6__ap_start;
  input Stream2Mmap_6__ap_ready;
  input Stream2Mmap_6__ap_done;
  input Stream2Mmap_6__ap_idle;
  output [63:0] Stream2Mmap_7___n__q0;
  output [63:0] Stream2Mmap_7___rmem7__q0;
  output Stream2Mmap_7__ap_start;
  input Stream2Mmap_7__ap_ready;
  input Stream2Mmap_7__ap_done;
  input Stream2Mmap_7__ap_idle;
  output [63:0] Stream2Mmap_8___n__q0;
  output [63:0] Stream2Mmap_8___rmem8__q0;
  output Stream2Mmap_8__ap_start;
  input Stream2Mmap_8__ap_ready;
  input Stream2Mmap_8__ap_done;
  input Stream2Mmap_8__ap_idle;
  output [63:0] Stream2Mmap_9___n__q0;
  output [63:0] Stream2Mmap_9___rmem9__q0;
  output Stream2Mmap_9__ap_start;
  input Stream2Mmap_9__ap_ready;
  input Stream2Mmap_9__ap_done;
  input Stream2Mmap_9__ap_idle;
  output [63:0] Stream2Mmap_10___n__q0;
  output [63:0] Stream2Mmap_10___rmem10__q0;
  output Stream2Mmap_10__ap_start;
  input Stream2Mmap_10__ap_ready;
  input Stream2Mmap_10__ap_done;
  input Stream2Mmap_10__ap_idle;
  output [63:0] Stream2Mmap_11___n__q0;
  output [63:0] Stream2Mmap_11___rmem11__q0;
  output Stream2Mmap_11__ap_start;
  input Stream2Mmap_11__ap_ready;
  input Stream2Mmap_11__ap_done;
  input Stream2Mmap_11__ap_idle;
  output [63:0] Stream2Mmap_12___n__q0;
  output [63:0] Stream2Mmap_12___rmem12__q0;
  output Stream2Mmap_12__ap_start;
  input Stream2Mmap_12__ap_ready;
  input Stream2Mmap_12__ap_done;
  input Stream2Mmap_12__ap_idle;
  output [63:0] Stream2Mmap_13___n__q0;
  output [63:0] Stream2Mmap_13___rmem13__q0;
  output Stream2Mmap_13__ap_start;
  input Stream2Mmap_13__ap_ready;
  input Stream2Mmap_13__ap_done;
  input Stream2Mmap_13__ap_idle;
  output [63:0] Stream2Mmap_14___n__q0;
  output [63:0] Stream2Mmap_14___rmem14__q0;
  output Stream2Mmap_14__ap_start;
  input Stream2Mmap_14__ap_ready;
  input Stream2Mmap_14__ap_done;
  input Stream2Mmap_14__ap_idle;
  output [63:0] Stream2Mmap_15___n__q0;
  output [63:0] Stream2Mmap_15___rmem15__q0;
  output Stream2Mmap_15__ap_start;
  input Stream2Mmap_15__ap_ready;
  input Stream2Mmap_15__ap_done;
  input Stream2Mmap_15__ap_idle;
  output [63:0] Stream2Mmap_16___n__q0;
  output [63:0] Stream2Mmap_16___rmem16__q0;
  output Stream2Mmap_16__ap_start;
  input Stream2Mmap_16__ap_ready;
  input Stream2Mmap_16__ap_done;
  input Stream2Mmap_16__ap_idle;
  output [63:0] Stream2Mmap_17___n__q0;
  output [63:0] Stream2Mmap_17___rmem17__q0;
  output Stream2Mmap_17__ap_start;
  input Stream2Mmap_17__ap_ready;
  input Stream2Mmap_17__ap_done;
  input Stream2Mmap_17__ap_idle;
  output [63:0] Stream2Mmap_18___n__q0;
  output [63:0] Stream2Mmap_18___rmem18__q0;
  output Stream2Mmap_18__ap_start;
  input Stream2Mmap_18__ap_ready;
  input Stream2Mmap_18__ap_done;
  input Stream2Mmap_18__ap_idle;
  output [63:0] Stream2Mmap_19___n__q0;
  output [63:0] Stream2Mmap_19___rmem19__q0;
  output Stream2Mmap_19__ap_start;
  input Stream2Mmap_19__ap_ready;
  input Stream2Mmap_19__ap_done;
  input Stream2Mmap_19__ap_idle;
  output [63:0] Stream2Mmap_20___n__q0;
  output [63:0] Stream2Mmap_20___rmem20__q0;
  output Stream2Mmap_20__ap_start;
  input Stream2Mmap_20__ap_ready;
  input Stream2Mmap_20__ap_done;
  input Stream2Mmap_20__ap_idle;
  output [63:0] Stream2Mmap_21___n__q0;
  output [63:0] Stream2Mmap_21___rmem21__q0;
  output Stream2Mmap_21__ap_start;
  input Stream2Mmap_21__ap_ready;
  input Stream2Mmap_21__ap_done;
  input Stream2Mmap_21__ap_idle;
  output [63:0] Stream2Mmap_22___n__q0;
  output [63:0] Stream2Mmap_22___rmem22__q0;
  output Stream2Mmap_22__ap_start;
  input Stream2Mmap_22__ap_ready;
  input Stream2Mmap_22__ap_done;
  input Stream2Mmap_22__ap_idle;
  output [63:0] Stream2Mmap_23___n__q0;
  output [63:0] Stream2Mmap_23___rmem23__q0;
  output Stream2Mmap_23__ap_start;
  input Stream2Mmap_23__ap_ready;
  input Stream2Mmap_23__ap_done;
  input Stream2Mmap_23__ap_idle;
  output [63:0] Stream2Mmap_24___n__q0;
  output [63:0] Stream2Mmap_24___rmem24__q0;
  output Stream2Mmap_24__ap_start;
  input Stream2Mmap_24__ap_ready;
  input Stream2Mmap_24__ap_done;
  input Stream2Mmap_24__ap_idle;
  output [63:0] Stream2Mmap_25___n__q0;
  output [63:0] Stream2Mmap_25___rmem25__q0;
  output Stream2Mmap_25__ap_start;
  input Stream2Mmap_25__ap_ready;
  input Stream2Mmap_25__ap_done;
  input Stream2Mmap_25__ap_idle;
  output [63:0] Stream2Mmap_26___n__q0;
  output [63:0] Stream2Mmap_26___rmem26__q0;
  output Stream2Mmap_26__ap_start;
  input Stream2Mmap_26__ap_ready;
  input Stream2Mmap_26__ap_done;
  input Stream2Mmap_26__ap_idle;
  output [63:0] yshift_0___n__q0;
  output yshift_0__ap_start;
  input yshift_0__ap_ready;
  input yshift_0__ap_done;
  input yshift_0__ap_idle;
  output [63:0] yshift_1___n__q0;
  output yshift_1__ap_start;
  input yshift_1__ap_ready;
  input yshift_1__ap_done;
  input yshift_1__ap_idle;
  output [63:0] yshift_2___n__q0;
  output yshift_2__ap_start;
  input yshift_2__ap_ready;
  input yshift_2__ap_done;
  input yshift_2__ap_idle;
  output [63:0] yshift_3___n__q0;
  output yshift_3__ap_start;
  input yshift_3__ap_ready;
  input yshift_3__ap_done;
  input yshift_3__ap_idle;
  output [63:0] yshift_4___n__q0;
  output yshift_4__ap_start;
  input yshift_4__ap_ready;
  input yshift_4__ap_done;
  input yshift_4__ap_idle;
  output [63:0] yshift_5___n__q0;
  output yshift_5__ap_start;
  input yshift_5__ap_ready;
  input yshift_5__ap_done;
  input yshift_5__ap_idle;
  output [63:0] yshift_6___n__q0;
  output yshift_6__ap_start;
  input yshift_6__ap_ready;
  input yshift_6__ap_done;
  input yshift_6__ap_idle;
  output [63:0] yshift_7___n__q0;
  output yshift_7__ap_start;
  input yshift_7__ap_ready;
  input yshift_7__ap_done;
  input yshift_7__ap_idle;
  output [63:0] yshift_8___n__q0;
  output yshift_8__ap_start;
  input yshift_8__ap_ready;
  input yshift_8__ap_done;
  input yshift_8__ap_idle;
  output [63:0] yshift_9___n__q0;
  output yshift_9__ap_start;
  input yshift_9__ap_ready;
  input yshift_9__ap_done;
  input yshift_9__ap_idle;
  output [63:0] yshift_10___n__q0;
  output yshift_10__ap_start;
  input yshift_10__ap_ready;
  input yshift_10__ap_done;
  input yshift_10__ap_idle;
  output [63:0] yshift_11___n__q0;
  output yshift_11__ap_start;
  input yshift_11__ap_ready;
  input yshift_11__ap_done;
  input yshift_11__ap_idle;
  output [63:0] yshift_12___n__q0;
  output yshift_12__ap_start;
  input yshift_12__ap_ready;
  input yshift_12__ap_done;
  input yshift_12__ap_idle;
  output [63:0] yshift_13___n__q0;
  output yshift_13__ap_start;
  input yshift_13__ap_ready;
  input yshift_13__ap_done;
  input yshift_13__ap_idle;
  output [63:0] yshift_14___n__q0;
  output yshift_14__ap_start;
  input yshift_14__ap_ready;
  input yshift_14__ap_done;
  input yshift_14__ap_idle;
  output [63:0] yshift_15___n__q0;
  output yshift_15__ap_start;
  input yshift_15__ap_ready;
  input yshift_15__ap_done;
  input yshift_15__ap_idle;
  output [63:0] yshift_16___n__q0;
  output yshift_16__ap_start;
  input yshift_16__ap_ready;
  input yshift_16__ap_done;
  input yshift_16__ap_idle;
  output [63:0] yshift_17___n__q0;
  output yshift_17__ap_start;
  input yshift_17__ap_ready;
  input yshift_17__ap_done;
  input yshift_17__ap_idle;
  output [63:0] yshift_18___n__q0;
  output yshift_18__ap_start;
  input yshift_18__ap_ready;
  input yshift_18__ap_done;
  input yshift_18__ap_idle;
  output [63:0] yshift_19___n__q0;
  output yshift_19__ap_start;
  input yshift_19__ap_ready;
  input yshift_19__ap_done;
  input yshift_19__ap_idle;
  output [63:0] yshift_20___n__q0;
  output yshift_20__ap_start;
  input yshift_20__ap_ready;
  input yshift_20__ap_done;
  input yshift_20__ap_idle;
  output [63:0] yshift_21___n__q0;
  output yshift_21__ap_start;
  input yshift_21__ap_ready;
  input yshift_21__ap_done;
  input yshift_21__ap_idle;
  output [63:0] yshift_22___n__q0;
  output yshift_22__ap_start;
  input yshift_22__ap_ready;
  input yshift_22__ap_done;
  input yshift_22__ap_idle;
  output [63:0] yshift_23___n__q0;
  output yshift_23__ap_start;
  input yshift_23__ap_ready;
  input yshift_23__ap_done;
  input yshift_23__ap_idle;
  output [63:0] yshift_24___n__q0;
  output yshift_24__ap_start;
  input yshift_24__ap_ready;
  input yshift_24__ap_done;
  input yshift_24__ap_idle;
  output [63:0] yshift_25___n__q0;
  output yshift_25__ap_start;
  input yshift_25__ap_ready;
  input yshift_25__ap_done;
  input yshift_25__ap_idle;
  output [63:0] yshift_26___n__q0;
  output yshift_26__ap_start;
  input yshift_26__ap_ready;
  input yshift_26__ap_done;
  input yshift_26__ap_idle;
  wire [63:0] Mmap2Stream_0___n__q0;
  wire [63:0] Mmap2Stream_0___rmem0__q0;
  wire Mmap2Stream_0__ap_start_global__q0;
  wire Mmap2Stream_0__is_done__q0;
  wire Mmap2Stream_0__ap_done_global__q0;
  wire Mmap2Stream_0__ap_start;
  wire Mmap2Stream_0__ap_ready;
  wire Mmap2Stream_0__ap_done;
  wire Mmap2Stream_0__ap_idle;
  reg [1:0] Mmap2Stream_0__state;
  wire [63:0] Mmap2Stream_1___n__q0;
  wire [63:0] Mmap2Stream_1___rmem1__q0;
  wire Mmap2Stream_1__ap_start_global__q0;
  wire Mmap2Stream_1__is_done__q0;
  wire Mmap2Stream_1__ap_done_global__q0;
  wire Mmap2Stream_1__ap_start;
  wire Mmap2Stream_1__ap_ready;
  wire Mmap2Stream_1__ap_done;
  wire Mmap2Stream_1__ap_idle;
  reg [1:0] Mmap2Stream_1__state;
  wire [63:0] Mmap2Stream_2___n__q0;
  wire [63:0] Mmap2Stream_2___rmem2__q0;
  wire Mmap2Stream_2__ap_start_global__q0;
  wire Mmap2Stream_2__is_done__q0;
  wire Mmap2Stream_2__ap_done_global__q0;
  wire Mmap2Stream_2__ap_start;
  wire Mmap2Stream_2__ap_ready;
  wire Mmap2Stream_2__ap_done;
  wire Mmap2Stream_2__ap_idle;
  reg [1:0] Mmap2Stream_2__state;
  wire [63:0] Mmap2Stream_3___n__q0;
  wire [63:0] Mmap2Stream_3___rmem3__q0;
  wire Mmap2Stream_3__ap_start_global__q0;
  wire Mmap2Stream_3__is_done__q0;
  wire Mmap2Stream_3__ap_done_global__q0;
  wire Mmap2Stream_3__ap_start;
  wire Mmap2Stream_3__ap_ready;
  wire Mmap2Stream_3__ap_done;
  wire Mmap2Stream_3__ap_idle;
  reg [1:0] Mmap2Stream_3__state;
  wire [63:0] Mmap2Stream_4___n__q0;
  wire [63:0] Mmap2Stream_4___rmem4__q0;
  wire Mmap2Stream_4__ap_start_global__q0;
  wire Mmap2Stream_4__is_done__q0;
  wire Mmap2Stream_4__ap_done_global__q0;
  wire Mmap2Stream_4__ap_start;
  wire Mmap2Stream_4__ap_ready;
  wire Mmap2Stream_4__ap_done;
  wire Mmap2Stream_4__ap_idle;
  reg [1:0] Mmap2Stream_4__state;
  wire [63:0] Mmap2Stream_5___n__q0;
  wire [63:0] Mmap2Stream_5___rmem5__q0;
  wire Mmap2Stream_5__ap_start_global__q0;
  wire Mmap2Stream_5__is_done__q0;
  wire Mmap2Stream_5__ap_done_global__q0;
  wire Mmap2Stream_5__ap_start;
  wire Mmap2Stream_5__ap_ready;
  wire Mmap2Stream_5__ap_done;
  wire Mmap2Stream_5__ap_idle;
  reg [1:0] Mmap2Stream_5__state;
  wire [63:0] Mmap2Stream_6___n__q0;
  wire [63:0] Mmap2Stream_6___rmem6__q0;
  wire Mmap2Stream_6__ap_start_global__q0;
  wire Mmap2Stream_6__is_done__q0;
  wire Mmap2Stream_6__ap_done_global__q0;
  wire Mmap2Stream_6__ap_start;
  wire Mmap2Stream_6__ap_ready;
  wire Mmap2Stream_6__ap_done;
  wire Mmap2Stream_6__ap_idle;
  reg [1:0] Mmap2Stream_6__state;
  wire [63:0] Mmap2Stream_7___n__q0;
  wire [63:0] Mmap2Stream_7___rmem7__q0;
  wire Mmap2Stream_7__ap_start_global__q0;
  wire Mmap2Stream_7__is_done__q0;
  wire Mmap2Stream_7__ap_done_global__q0;
  wire Mmap2Stream_7__ap_start;
  wire Mmap2Stream_7__ap_ready;
  wire Mmap2Stream_7__ap_done;
  wire Mmap2Stream_7__ap_idle;
  reg [1:0] Mmap2Stream_7__state;
  wire [63:0] Mmap2Stream_8___n__q0;
  wire [63:0] Mmap2Stream_8___rmem8__q0;
  wire Mmap2Stream_8__ap_start_global__q0;
  wire Mmap2Stream_8__is_done__q0;
  wire Mmap2Stream_8__ap_done_global__q0;
  wire Mmap2Stream_8__ap_start;
  wire Mmap2Stream_8__ap_ready;
  wire Mmap2Stream_8__ap_done;
  wire Mmap2Stream_8__ap_idle;
  reg [1:0] Mmap2Stream_8__state;
  wire [63:0] Mmap2Stream_9___n__q0;
  wire [63:0] Mmap2Stream_9___rmem9__q0;
  wire Mmap2Stream_9__ap_start_global__q0;
  wire Mmap2Stream_9__is_done__q0;
  wire Mmap2Stream_9__ap_done_global__q0;
  wire Mmap2Stream_9__ap_start;
  wire Mmap2Stream_9__ap_ready;
  wire Mmap2Stream_9__ap_done;
  wire Mmap2Stream_9__ap_idle;
  reg [1:0] Mmap2Stream_9__state;
  wire [63:0] Mmap2Stream_10___n__q0;
  wire [63:0] Mmap2Stream_10___rmem10__q0;
  wire Mmap2Stream_10__ap_start_global__q0;
  wire Mmap2Stream_10__is_done__q0;
  wire Mmap2Stream_10__ap_done_global__q0;
  wire Mmap2Stream_10__ap_start;
  wire Mmap2Stream_10__ap_ready;
  wire Mmap2Stream_10__ap_done;
  wire Mmap2Stream_10__ap_idle;
  reg [1:0] Mmap2Stream_10__state;
  wire [63:0] Mmap2Stream_11___n__q0;
  wire [63:0] Mmap2Stream_11___rmem11__q0;
  wire Mmap2Stream_11__ap_start_global__q0;
  wire Mmap2Stream_11__is_done__q0;
  wire Mmap2Stream_11__ap_done_global__q0;
  wire Mmap2Stream_11__ap_start;
  wire Mmap2Stream_11__ap_ready;
  wire Mmap2Stream_11__ap_done;
  wire Mmap2Stream_11__ap_idle;
  reg [1:0] Mmap2Stream_11__state;
  wire [63:0] Mmap2Stream_12___n__q0;
  wire [63:0] Mmap2Stream_12___rmem12__q0;
  wire Mmap2Stream_12__ap_start_global__q0;
  wire Mmap2Stream_12__is_done__q0;
  wire Mmap2Stream_12__ap_done_global__q0;
  wire Mmap2Stream_12__ap_start;
  wire Mmap2Stream_12__ap_ready;
  wire Mmap2Stream_12__ap_done;
  wire Mmap2Stream_12__ap_idle;
  reg [1:0] Mmap2Stream_12__state;
  wire [63:0] Mmap2Stream_13___n__q0;
  wire [63:0] Mmap2Stream_13___rmem13__q0;
  wire Mmap2Stream_13__ap_start_global__q0;
  wire Mmap2Stream_13__is_done__q0;
  wire Mmap2Stream_13__ap_done_global__q0;
  wire Mmap2Stream_13__ap_start;
  wire Mmap2Stream_13__ap_ready;
  wire Mmap2Stream_13__ap_done;
  wire Mmap2Stream_13__ap_idle;
  reg [1:0] Mmap2Stream_13__state;
  wire [63:0] Mmap2Stream_14___n__q0;
  wire [63:0] Mmap2Stream_14___rmem14__q0;
  wire Mmap2Stream_14__ap_start_global__q0;
  wire Mmap2Stream_14__is_done__q0;
  wire Mmap2Stream_14__ap_done_global__q0;
  wire Mmap2Stream_14__ap_start;
  wire Mmap2Stream_14__ap_ready;
  wire Mmap2Stream_14__ap_done;
  wire Mmap2Stream_14__ap_idle;
  reg [1:0] Mmap2Stream_14__state;
  wire [63:0] Mmap2Stream_15___n__q0;
  wire [63:0] Mmap2Stream_15___rmem15__q0;
  wire Mmap2Stream_15__ap_start_global__q0;
  wire Mmap2Stream_15__is_done__q0;
  wire Mmap2Stream_15__ap_done_global__q0;
  wire Mmap2Stream_15__ap_start;
  wire Mmap2Stream_15__ap_ready;
  wire Mmap2Stream_15__ap_done;
  wire Mmap2Stream_15__ap_idle;
  reg [1:0] Mmap2Stream_15__state;
  wire [63:0] Mmap2Stream_16___n__q0;
  wire [63:0] Mmap2Stream_16___rmem16__q0;
  wire Mmap2Stream_16__ap_start_global__q0;
  wire Mmap2Stream_16__is_done__q0;
  wire Mmap2Stream_16__ap_done_global__q0;
  wire Mmap2Stream_16__ap_start;
  wire Mmap2Stream_16__ap_ready;
  wire Mmap2Stream_16__ap_done;
  wire Mmap2Stream_16__ap_idle;
  reg [1:0] Mmap2Stream_16__state;
  wire [63:0] Mmap2Stream_17___n__q0;
  wire [63:0] Mmap2Stream_17___rmem17__q0;
  wire Mmap2Stream_17__ap_start_global__q0;
  wire Mmap2Stream_17__is_done__q0;
  wire Mmap2Stream_17__ap_done_global__q0;
  wire Mmap2Stream_17__ap_start;
  wire Mmap2Stream_17__ap_ready;
  wire Mmap2Stream_17__ap_done;
  wire Mmap2Stream_17__ap_idle;
  reg [1:0] Mmap2Stream_17__state;
  wire [63:0] Mmap2Stream_18___n__q0;
  wire [63:0] Mmap2Stream_18___rmem18__q0;
  wire Mmap2Stream_18__ap_start_global__q0;
  wire Mmap2Stream_18__is_done__q0;
  wire Mmap2Stream_18__ap_done_global__q0;
  wire Mmap2Stream_18__ap_start;
  wire Mmap2Stream_18__ap_ready;
  wire Mmap2Stream_18__ap_done;
  wire Mmap2Stream_18__ap_idle;
  reg [1:0] Mmap2Stream_18__state;
  wire [63:0] Mmap2Stream_19___n__q0;
  wire [63:0] Mmap2Stream_19___rmem19__q0;
  wire Mmap2Stream_19__ap_start_global__q0;
  wire Mmap2Stream_19__is_done__q0;
  wire Mmap2Stream_19__ap_done_global__q0;
  wire Mmap2Stream_19__ap_start;
  wire Mmap2Stream_19__ap_ready;
  wire Mmap2Stream_19__ap_done;
  wire Mmap2Stream_19__ap_idle;
  reg [1:0] Mmap2Stream_19__state;
  wire [63:0] Mmap2Stream_20___n__q0;
  wire [63:0] Mmap2Stream_20___rmem20__q0;
  wire Mmap2Stream_20__ap_start_global__q0;
  wire Mmap2Stream_20__is_done__q0;
  wire Mmap2Stream_20__ap_done_global__q0;
  wire Mmap2Stream_20__ap_start;
  wire Mmap2Stream_20__ap_ready;
  wire Mmap2Stream_20__ap_done;
  wire Mmap2Stream_20__ap_idle;
  reg [1:0] Mmap2Stream_20__state;
  wire [63:0] Mmap2Stream_21___n__q0;
  wire [63:0] Mmap2Stream_21___rmem21__q0;
  wire Mmap2Stream_21__ap_start_global__q0;
  wire Mmap2Stream_21__is_done__q0;
  wire Mmap2Stream_21__ap_done_global__q0;
  wire Mmap2Stream_21__ap_start;
  wire Mmap2Stream_21__ap_ready;
  wire Mmap2Stream_21__ap_done;
  wire Mmap2Stream_21__ap_idle;
  reg [1:0] Mmap2Stream_21__state;
  wire [63:0] Mmap2Stream_22___n__q0;
  wire [63:0] Mmap2Stream_22___rmem22__q0;
  wire Mmap2Stream_22__ap_start_global__q0;
  wire Mmap2Stream_22__is_done__q0;
  wire Mmap2Stream_22__ap_done_global__q0;
  wire Mmap2Stream_22__ap_start;
  wire Mmap2Stream_22__ap_ready;
  wire Mmap2Stream_22__ap_done;
  wire Mmap2Stream_22__ap_idle;
  reg [1:0] Mmap2Stream_22__state;
  wire [63:0] Mmap2Stream_23___n__q0;
  wire [63:0] Mmap2Stream_23___rmem23__q0;
  wire Mmap2Stream_23__ap_start_global__q0;
  wire Mmap2Stream_23__is_done__q0;
  wire Mmap2Stream_23__ap_done_global__q0;
  wire Mmap2Stream_23__ap_start;
  wire Mmap2Stream_23__ap_ready;
  wire Mmap2Stream_23__ap_done;
  wire Mmap2Stream_23__ap_idle;
  reg [1:0] Mmap2Stream_23__state;
  wire [63:0] Mmap2Stream_24___n__q0;
  wire [63:0] Mmap2Stream_24___rmem24__q0;
  wire Mmap2Stream_24__ap_start_global__q0;
  wire Mmap2Stream_24__is_done__q0;
  wire Mmap2Stream_24__ap_done_global__q0;
  wire Mmap2Stream_24__ap_start;
  wire Mmap2Stream_24__ap_ready;
  wire Mmap2Stream_24__ap_done;
  wire Mmap2Stream_24__ap_idle;
  reg [1:0] Mmap2Stream_24__state;
  wire [63:0] Mmap2Stream_25___n__q0;
  wire [63:0] Mmap2Stream_25___rmem25__q0;
  wire Mmap2Stream_25__ap_start_global__q0;
  wire Mmap2Stream_25__is_done__q0;
  wire Mmap2Stream_25__ap_done_global__q0;
  wire Mmap2Stream_25__ap_start;
  wire Mmap2Stream_25__ap_ready;
  wire Mmap2Stream_25__ap_done;
  wire Mmap2Stream_25__ap_idle;
  reg [1:0] Mmap2Stream_25__state;
  wire [63:0] Mmap2Stream_26___n__q0;
  wire [63:0] Mmap2Stream_26___rmem26__q0;
  wire Mmap2Stream_26__ap_start_global__q0;
  wire Mmap2Stream_26__is_done__q0;
  wire Mmap2Stream_26__ap_done_global__q0;
  wire Mmap2Stream_26__ap_start;
  wire Mmap2Stream_26__ap_ready;
  wire Mmap2Stream_26__ap_done;
  wire Mmap2Stream_26__ap_idle;
  reg [1:0] Mmap2Stream_26__state;
  wire [63:0] Stream2Mmap_0___n__q0;
  wire [63:0] Stream2Mmap_0___rmem0__q0;
  wire Stream2Mmap_0__ap_start_global__q0;
  wire Stream2Mmap_0__is_done__q0;
  wire Stream2Mmap_0__ap_done_global__q0;
  wire Stream2Mmap_0__ap_start;
  wire Stream2Mmap_0__ap_ready;
  wire Stream2Mmap_0__ap_done;
  wire Stream2Mmap_0__ap_idle;
  reg [1:0] Stream2Mmap_0__state;
  wire [63:0] Stream2Mmap_1___n__q0;
  wire [63:0] Stream2Mmap_1___rmem1__q0;
  wire Stream2Mmap_1__ap_start_global__q0;
  wire Stream2Mmap_1__is_done__q0;
  wire Stream2Mmap_1__ap_done_global__q0;
  wire Stream2Mmap_1__ap_start;
  wire Stream2Mmap_1__ap_ready;
  wire Stream2Mmap_1__ap_done;
  wire Stream2Mmap_1__ap_idle;
  reg [1:0] Stream2Mmap_1__state;
  wire [63:0] Stream2Mmap_2___n__q0;
  wire [63:0] Stream2Mmap_2___rmem2__q0;
  wire Stream2Mmap_2__ap_start_global__q0;
  wire Stream2Mmap_2__is_done__q0;
  wire Stream2Mmap_2__ap_done_global__q0;
  wire Stream2Mmap_2__ap_start;
  wire Stream2Mmap_2__ap_ready;
  wire Stream2Mmap_2__ap_done;
  wire Stream2Mmap_2__ap_idle;
  reg [1:0] Stream2Mmap_2__state;
  wire [63:0] Stream2Mmap_3___n__q0;
  wire [63:0] Stream2Mmap_3___rmem3__q0;
  wire Stream2Mmap_3__ap_start_global__q0;
  wire Stream2Mmap_3__is_done__q0;
  wire Stream2Mmap_3__ap_done_global__q0;
  wire Stream2Mmap_3__ap_start;
  wire Stream2Mmap_3__ap_ready;
  wire Stream2Mmap_3__ap_done;
  wire Stream2Mmap_3__ap_idle;
  reg [1:0] Stream2Mmap_3__state;
  wire [63:0] Stream2Mmap_4___n__q0;
  wire [63:0] Stream2Mmap_4___rmem4__q0;
  wire Stream2Mmap_4__ap_start_global__q0;
  wire Stream2Mmap_4__is_done__q0;
  wire Stream2Mmap_4__ap_done_global__q0;
  wire Stream2Mmap_4__ap_start;
  wire Stream2Mmap_4__ap_ready;
  wire Stream2Mmap_4__ap_done;
  wire Stream2Mmap_4__ap_idle;
  reg [1:0] Stream2Mmap_4__state;
  wire [63:0] Stream2Mmap_5___n__q0;
  wire [63:0] Stream2Mmap_5___rmem5__q0;
  wire Stream2Mmap_5__ap_start_global__q0;
  wire Stream2Mmap_5__is_done__q0;
  wire Stream2Mmap_5__ap_done_global__q0;
  wire Stream2Mmap_5__ap_start;
  wire Stream2Mmap_5__ap_ready;
  wire Stream2Mmap_5__ap_done;
  wire Stream2Mmap_5__ap_idle;
  reg [1:0] Stream2Mmap_5__state;
  wire [63:0] Stream2Mmap_6___n__q0;
  wire [63:0] Stream2Mmap_6___rmem6__q0;
  wire Stream2Mmap_6__ap_start_global__q0;
  wire Stream2Mmap_6__is_done__q0;
  wire Stream2Mmap_6__ap_done_global__q0;
  wire Stream2Mmap_6__ap_start;
  wire Stream2Mmap_6__ap_ready;
  wire Stream2Mmap_6__ap_done;
  wire Stream2Mmap_6__ap_idle;
  reg [1:0] Stream2Mmap_6__state;
  wire [63:0] Stream2Mmap_7___n__q0;
  wire [63:0] Stream2Mmap_7___rmem7__q0;
  wire Stream2Mmap_7__ap_start_global__q0;
  wire Stream2Mmap_7__is_done__q0;
  wire Stream2Mmap_7__ap_done_global__q0;
  wire Stream2Mmap_7__ap_start;
  wire Stream2Mmap_7__ap_ready;
  wire Stream2Mmap_7__ap_done;
  wire Stream2Mmap_7__ap_idle;
  reg [1:0] Stream2Mmap_7__state;
  wire [63:0] Stream2Mmap_8___n__q0;
  wire [63:0] Stream2Mmap_8___rmem8__q0;
  wire Stream2Mmap_8__ap_start_global__q0;
  wire Stream2Mmap_8__is_done__q0;
  wire Stream2Mmap_8__ap_done_global__q0;
  wire Stream2Mmap_8__ap_start;
  wire Stream2Mmap_8__ap_ready;
  wire Stream2Mmap_8__ap_done;
  wire Stream2Mmap_8__ap_idle;
  reg [1:0] Stream2Mmap_8__state;
  wire [63:0] Stream2Mmap_9___n__q0;
  wire [63:0] Stream2Mmap_9___rmem9__q0;
  wire Stream2Mmap_9__ap_start_global__q0;
  wire Stream2Mmap_9__is_done__q0;
  wire Stream2Mmap_9__ap_done_global__q0;
  wire Stream2Mmap_9__ap_start;
  wire Stream2Mmap_9__ap_ready;
  wire Stream2Mmap_9__ap_done;
  wire Stream2Mmap_9__ap_idle;
  reg [1:0] Stream2Mmap_9__state;
  wire [63:0] Stream2Mmap_10___n__q0;
  wire [63:0] Stream2Mmap_10___rmem10__q0;
  wire Stream2Mmap_10__ap_start_global__q0;
  wire Stream2Mmap_10__is_done__q0;
  wire Stream2Mmap_10__ap_done_global__q0;
  wire Stream2Mmap_10__ap_start;
  wire Stream2Mmap_10__ap_ready;
  wire Stream2Mmap_10__ap_done;
  wire Stream2Mmap_10__ap_idle;
  reg [1:0] Stream2Mmap_10__state;
  wire [63:0] Stream2Mmap_11___n__q0;
  wire [63:0] Stream2Mmap_11___rmem11__q0;
  wire Stream2Mmap_11__ap_start_global__q0;
  wire Stream2Mmap_11__is_done__q0;
  wire Stream2Mmap_11__ap_done_global__q0;
  wire Stream2Mmap_11__ap_start;
  wire Stream2Mmap_11__ap_ready;
  wire Stream2Mmap_11__ap_done;
  wire Stream2Mmap_11__ap_idle;
  reg [1:0] Stream2Mmap_11__state;
  wire [63:0] Stream2Mmap_12___n__q0;
  wire [63:0] Stream2Mmap_12___rmem12__q0;
  wire Stream2Mmap_12__ap_start_global__q0;
  wire Stream2Mmap_12__is_done__q0;
  wire Stream2Mmap_12__ap_done_global__q0;
  wire Stream2Mmap_12__ap_start;
  wire Stream2Mmap_12__ap_ready;
  wire Stream2Mmap_12__ap_done;
  wire Stream2Mmap_12__ap_idle;
  reg [1:0] Stream2Mmap_12__state;
  wire [63:0] Stream2Mmap_13___n__q0;
  wire [63:0] Stream2Mmap_13___rmem13__q0;
  wire Stream2Mmap_13__ap_start_global__q0;
  wire Stream2Mmap_13__is_done__q0;
  wire Stream2Mmap_13__ap_done_global__q0;
  wire Stream2Mmap_13__ap_start;
  wire Stream2Mmap_13__ap_ready;
  wire Stream2Mmap_13__ap_done;
  wire Stream2Mmap_13__ap_idle;
  reg [1:0] Stream2Mmap_13__state;
  wire [63:0] Stream2Mmap_14___n__q0;
  wire [63:0] Stream2Mmap_14___rmem14__q0;
  wire Stream2Mmap_14__ap_start_global__q0;
  wire Stream2Mmap_14__is_done__q0;
  wire Stream2Mmap_14__ap_done_global__q0;
  wire Stream2Mmap_14__ap_start;
  wire Stream2Mmap_14__ap_ready;
  wire Stream2Mmap_14__ap_done;
  wire Stream2Mmap_14__ap_idle;
  reg [1:0] Stream2Mmap_14__state;
  wire [63:0] Stream2Mmap_15___n__q0;
  wire [63:0] Stream2Mmap_15___rmem15__q0;
  wire Stream2Mmap_15__ap_start_global__q0;
  wire Stream2Mmap_15__is_done__q0;
  wire Stream2Mmap_15__ap_done_global__q0;
  wire Stream2Mmap_15__ap_start;
  wire Stream2Mmap_15__ap_ready;
  wire Stream2Mmap_15__ap_done;
  wire Stream2Mmap_15__ap_idle;
  reg [1:0] Stream2Mmap_15__state;
  wire [63:0] Stream2Mmap_16___n__q0;
  wire [63:0] Stream2Mmap_16___rmem16__q0;
  wire Stream2Mmap_16__ap_start_global__q0;
  wire Stream2Mmap_16__is_done__q0;
  wire Stream2Mmap_16__ap_done_global__q0;
  wire Stream2Mmap_16__ap_start;
  wire Stream2Mmap_16__ap_ready;
  wire Stream2Mmap_16__ap_done;
  wire Stream2Mmap_16__ap_idle;
  reg [1:0] Stream2Mmap_16__state;
  wire [63:0] Stream2Mmap_17___n__q0;
  wire [63:0] Stream2Mmap_17___rmem17__q0;
  wire Stream2Mmap_17__ap_start_global__q0;
  wire Stream2Mmap_17__is_done__q0;
  wire Stream2Mmap_17__ap_done_global__q0;
  wire Stream2Mmap_17__ap_start;
  wire Stream2Mmap_17__ap_ready;
  wire Stream2Mmap_17__ap_done;
  wire Stream2Mmap_17__ap_idle;
  reg [1:0] Stream2Mmap_17__state;
  wire [63:0] Stream2Mmap_18___n__q0;
  wire [63:0] Stream2Mmap_18___rmem18__q0;
  wire Stream2Mmap_18__ap_start_global__q0;
  wire Stream2Mmap_18__is_done__q0;
  wire Stream2Mmap_18__ap_done_global__q0;
  wire Stream2Mmap_18__ap_start;
  wire Stream2Mmap_18__ap_ready;
  wire Stream2Mmap_18__ap_done;
  wire Stream2Mmap_18__ap_idle;
  reg [1:0] Stream2Mmap_18__state;
  wire [63:0] Stream2Mmap_19___n__q0;
  wire [63:0] Stream2Mmap_19___rmem19__q0;
  wire Stream2Mmap_19__ap_start_global__q0;
  wire Stream2Mmap_19__is_done__q0;
  wire Stream2Mmap_19__ap_done_global__q0;
  wire Stream2Mmap_19__ap_start;
  wire Stream2Mmap_19__ap_ready;
  wire Stream2Mmap_19__ap_done;
  wire Stream2Mmap_19__ap_idle;
  reg [1:0] Stream2Mmap_19__state;
  wire [63:0] Stream2Mmap_20___n__q0;
  wire [63:0] Stream2Mmap_20___rmem20__q0;
  wire Stream2Mmap_20__ap_start_global__q0;
  wire Stream2Mmap_20__is_done__q0;
  wire Stream2Mmap_20__ap_done_global__q0;
  wire Stream2Mmap_20__ap_start;
  wire Stream2Mmap_20__ap_ready;
  wire Stream2Mmap_20__ap_done;
  wire Stream2Mmap_20__ap_idle;
  reg [1:0] Stream2Mmap_20__state;
  wire [63:0] Stream2Mmap_21___n__q0;
  wire [63:0] Stream2Mmap_21___rmem21__q0;
  wire Stream2Mmap_21__ap_start_global__q0;
  wire Stream2Mmap_21__is_done__q0;
  wire Stream2Mmap_21__ap_done_global__q0;
  wire Stream2Mmap_21__ap_start;
  wire Stream2Mmap_21__ap_ready;
  wire Stream2Mmap_21__ap_done;
  wire Stream2Mmap_21__ap_idle;
  reg [1:0] Stream2Mmap_21__state;
  wire [63:0] Stream2Mmap_22___n__q0;
  wire [63:0] Stream2Mmap_22___rmem22__q0;
  wire Stream2Mmap_22__ap_start_global__q0;
  wire Stream2Mmap_22__is_done__q0;
  wire Stream2Mmap_22__ap_done_global__q0;
  wire Stream2Mmap_22__ap_start;
  wire Stream2Mmap_22__ap_ready;
  wire Stream2Mmap_22__ap_done;
  wire Stream2Mmap_22__ap_idle;
  reg [1:0] Stream2Mmap_22__state;
  wire [63:0] Stream2Mmap_23___n__q0;
  wire [63:0] Stream2Mmap_23___rmem23__q0;
  wire Stream2Mmap_23__ap_start_global__q0;
  wire Stream2Mmap_23__is_done__q0;
  wire Stream2Mmap_23__ap_done_global__q0;
  wire Stream2Mmap_23__ap_start;
  wire Stream2Mmap_23__ap_ready;
  wire Stream2Mmap_23__ap_done;
  wire Stream2Mmap_23__ap_idle;
  reg [1:0] Stream2Mmap_23__state;
  wire [63:0] Stream2Mmap_24___n__q0;
  wire [63:0] Stream2Mmap_24___rmem24__q0;
  wire Stream2Mmap_24__ap_start_global__q0;
  wire Stream2Mmap_24__is_done__q0;
  wire Stream2Mmap_24__ap_done_global__q0;
  wire Stream2Mmap_24__ap_start;
  wire Stream2Mmap_24__ap_ready;
  wire Stream2Mmap_24__ap_done;
  wire Stream2Mmap_24__ap_idle;
  reg [1:0] Stream2Mmap_24__state;
  wire [63:0] Stream2Mmap_25___n__q0;
  wire [63:0] Stream2Mmap_25___rmem25__q0;
  wire Stream2Mmap_25__ap_start_global__q0;
  wire Stream2Mmap_25__is_done__q0;
  wire Stream2Mmap_25__ap_done_global__q0;
  wire Stream2Mmap_25__ap_start;
  wire Stream2Mmap_25__ap_ready;
  wire Stream2Mmap_25__ap_done;
  wire Stream2Mmap_25__ap_idle;
  reg [1:0] Stream2Mmap_25__state;
  wire [63:0] Stream2Mmap_26___n__q0;
  wire [63:0] Stream2Mmap_26___rmem26__q0;
  wire Stream2Mmap_26__ap_start_global__q0;
  wire Stream2Mmap_26__is_done__q0;
  wire Stream2Mmap_26__ap_done_global__q0;
  wire Stream2Mmap_26__ap_start;
  wire Stream2Mmap_26__ap_ready;
  wire Stream2Mmap_26__ap_done;
  wire Stream2Mmap_26__ap_idle;
  reg [1:0] Stream2Mmap_26__state;
  wire [63:0] yshift_0___n__q0;
  wire yshift_0__ap_start_global__q0;
  wire yshift_0__is_done__q0;
  wire yshift_0__ap_done_global__q0;
  wire yshift_0__ap_start;
  wire yshift_0__ap_ready;
  wire yshift_0__ap_done;
  wire yshift_0__ap_idle;
  reg [1:0] yshift_0__state;
  wire [63:0] yshift_1___n__q0;
  wire yshift_1__ap_start_global__q0;
  wire yshift_1__is_done__q0;
  wire yshift_1__ap_done_global__q0;
  wire yshift_1__ap_start;
  wire yshift_1__ap_ready;
  wire yshift_1__ap_done;
  wire yshift_1__ap_idle;
  reg [1:0] yshift_1__state;
  wire [63:0] yshift_2___n__q0;
  wire yshift_2__ap_start_global__q0;
  wire yshift_2__is_done__q0;
  wire yshift_2__ap_done_global__q0;
  wire yshift_2__ap_start;
  wire yshift_2__ap_ready;
  wire yshift_2__ap_done;
  wire yshift_2__ap_idle;
  reg [1:0] yshift_2__state;
  wire [63:0] yshift_3___n__q0;
  wire yshift_3__ap_start_global__q0;
  wire yshift_3__is_done__q0;
  wire yshift_3__ap_done_global__q0;
  wire yshift_3__ap_start;
  wire yshift_3__ap_ready;
  wire yshift_3__ap_done;
  wire yshift_3__ap_idle;
  reg [1:0] yshift_3__state;
  wire [63:0] yshift_4___n__q0;
  wire yshift_4__ap_start_global__q0;
  wire yshift_4__is_done__q0;
  wire yshift_4__ap_done_global__q0;
  wire yshift_4__ap_start;
  wire yshift_4__ap_ready;
  wire yshift_4__ap_done;
  wire yshift_4__ap_idle;
  reg [1:0] yshift_4__state;
  wire [63:0] yshift_5___n__q0;
  wire yshift_5__ap_start_global__q0;
  wire yshift_5__is_done__q0;
  wire yshift_5__ap_done_global__q0;
  wire yshift_5__ap_start;
  wire yshift_5__ap_ready;
  wire yshift_5__ap_done;
  wire yshift_5__ap_idle;
  reg [1:0] yshift_5__state;
  wire [63:0] yshift_6___n__q0;
  wire yshift_6__ap_start_global__q0;
  wire yshift_6__is_done__q0;
  wire yshift_6__ap_done_global__q0;
  wire yshift_6__ap_start;
  wire yshift_6__ap_ready;
  wire yshift_6__ap_done;
  wire yshift_6__ap_idle;
  reg [1:0] yshift_6__state;
  wire [63:0] yshift_7___n__q0;
  wire yshift_7__ap_start_global__q0;
  wire yshift_7__is_done__q0;
  wire yshift_7__ap_done_global__q0;
  wire yshift_7__ap_start;
  wire yshift_7__ap_ready;
  wire yshift_7__ap_done;
  wire yshift_7__ap_idle;
  reg [1:0] yshift_7__state;
  wire [63:0] yshift_8___n__q0;
  wire yshift_8__ap_start_global__q0;
  wire yshift_8__is_done__q0;
  wire yshift_8__ap_done_global__q0;
  wire yshift_8__ap_start;
  wire yshift_8__ap_ready;
  wire yshift_8__ap_done;
  wire yshift_8__ap_idle;
  reg [1:0] yshift_8__state;
  wire [63:0] yshift_9___n__q0;
  wire yshift_9__ap_start_global__q0;
  wire yshift_9__is_done__q0;
  wire yshift_9__ap_done_global__q0;
  wire yshift_9__ap_start;
  wire yshift_9__ap_ready;
  wire yshift_9__ap_done;
  wire yshift_9__ap_idle;
  reg [1:0] yshift_9__state;
  wire [63:0] yshift_10___n__q0;
  wire yshift_10__ap_start_global__q0;
  wire yshift_10__is_done__q0;
  wire yshift_10__ap_done_global__q0;
  wire yshift_10__ap_start;
  wire yshift_10__ap_ready;
  wire yshift_10__ap_done;
  wire yshift_10__ap_idle;
  reg [1:0] yshift_10__state;
  wire [63:0] yshift_11___n__q0;
  wire yshift_11__ap_start_global__q0;
  wire yshift_11__is_done__q0;
  wire yshift_11__ap_done_global__q0;
  wire yshift_11__ap_start;
  wire yshift_11__ap_ready;
  wire yshift_11__ap_done;
  wire yshift_11__ap_idle;
  reg [1:0] yshift_11__state;
  wire [63:0] yshift_12___n__q0;
  wire yshift_12__ap_start_global__q0;
  wire yshift_12__is_done__q0;
  wire yshift_12__ap_done_global__q0;
  wire yshift_12__ap_start;
  wire yshift_12__ap_ready;
  wire yshift_12__ap_done;
  wire yshift_12__ap_idle;
  reg [1:0] yshift_12__state;
  wire [63:0] yshift_13___n__q0;
  wire yshift_13__ap_start_global__q0;
  wire yshift_13__is_done__q0;
  wire yshift_13__ap_done_global__q0;
  wire yshift_13__ap_start;
  wire yshift_13__ap_ready;
  wire yshift_13__ap_done;
  wire yshift_13__ap_idle;
  reg [1:0] yshift_13__state;
  wire [63:0] yshift_14___n__q0;
  wire yshift_14__ap_start_global__q0;
  wire yshift_14__is_done__q0;
  wire yshift_14__ap_done_global__q0;
  wire yshift_14__ap_start;
  wire yshift_14__ap_ready;
  wire yshift_14__ap_done;
  wire yshift_14__ap_idle;
  reg [1:0] yshift_14__state;
  wire [63:0] yshift_15___n__q0;
  wire yshift_15__ap_start_global__q0;
  wire yshift_15__is_done__q0;
  wire yshift_15__ap_done_global__q0;
  wire yshift_15__ap_start;
  wire yshift_15__ap_ready;
  wire yshift_15__ap_done;
  wire yshift_15__ap_idle;
  reg [1:0] yshift_15__state;
  wire [63:0] yshift_16___n__q0;
  wire yshift_16__ap_start_global__q0;
  wire yshift_16__is_done__q0;
  wire yshift_16__ap_done_global__q0;
  wire yshift_16__ap_start;
  wire yshift_16__ap_ready;
  wire yshift_16__ap_done;
  wire yshift_16__ap_idle;
  reg [1:0] yshift_16__state;
  wire [63:0] yshift_17___n__q0;
  wire yshift_17__ap_start_global__q0;
  wire yshift_17__is_done__q0;
  wire yshift_17__ap_done_global__q0;
  wire yshift_17__ap_start;
  wire yshift_17__ap_ready;
  wire yshift_17__ap_done;
  wire yshift_17__ap_idle;
  reg [1:0] yshift_17__state;
  wire [63:0] yshift_18___n__q0;
  wire yshift_18__ap_start_global__q0;
  wire yshift_18__is_done__q0;
  wire yshift_18__ap_done_global__q0;
  wire yshift_18__ap_start;
  wire yshift_18__ap_ready;
  wire yshift_18__ap_done;
  wire yshift_18__ap_idle;
  reg [1:0] yshift_18__state;
  wire [63:0] yshift_19___n__q0;
  wire yshift_19__ap_start_global__q0;
  wire yshift_19__is_done__q0;
  wire yshift_19__ap_done_global__q0;
  wire yshift_19__ap_start;
  wire yshift_19__ap_ready;
  wire yshift_19__ap_done;
  wire yshift_19__ap_idle;
  reg [1:0] yshift_19__state;
  wire [63:0] yshift_20___n__q0;
  wire yshift_20__ap_start_global__q0;
  wire yshift_20__is_done__q0;
  wire yshift_20__ap_done_global__q0;
  wire yshift_20__ap_start;
  wire yshift_20__ap_ready;
  wire yshift_20__ap_done;
  wire yshift_20__ap_idle;
  reg [1:0] yshift_20__state;
  wire [63:0] yshift_21___n__q0;
  wire yshift_21__ap_start_global__q0;
  wire yshift_21__is_done__q0;
  wire yshift_21__ap_done_global__q0;
  wire yshift_21__ap_start;
  wire yshift_21__ap_ready;
  wire yshift_21__ap_done;
  wire yshift_21__ap_idle;
  reg [1:0] yshift_21__state;
  wire [63:0] yshift_22___n__q0;
  wire yshift_22__ap_start_global__q0;
  wire yshift_22__is_done__q0;
  wire yshift_22__ap_done_global__q0;
  wire yshift_22__ap_start;
  wire yshift_22__ap_ready;
  wire yshift_22__ap_done;
  wire yshift_22__ap_idle;
  reg [1:0] yshift_22__state;
  wire [63:0] yshift_23___n__q0;
  wire yshift_23__ap_start_global__q0;
  wire yshift_23__is_done__q0;
  wire yshift_23__ap_done_global__q0;
  wire yshift_23__ap_start;
  wire yshift_23__ap_ready;
  wire yshift_23__ap_done;
  wire yshift_23__ap_idle;
  reg [1:0] yshift_23__state;
  wire [63:0] yshift_24___n__q0;
  wire yshift_24__ap_start_global__q0;
  wire yshift_24__is_done__q0;
  wire yshift_24__ap_done_global__q0;
  wire yshift_24__ap_start;
  wire yshift_24__ap_ready;
  wire yshift_24__ap_done;
  wire yshift_24__ap_idle;
  reg [1:0] yshift_24__state;
  wire [63:0] yshift_25___n__q0;
  wire yshift_25__ap_start_global__q0;
  wire yshift_25__is_done__q0;
  wire yshift_25__ap_done_global__q0;
  wire yshift_25__ap_start;
  wire yshift_25__ap_ready;
  wire yshift_25__ap_done;
  wire yshift_25__ap_idle;
  reg [1:0] yshift_25__state;
  wire [63:0] yshift_26___n__q0;
  wire yshift_26__ap_start_global__q0;
  wire yshift_26__is_done__q0;
  wire yshift_26__ap_done_global__q0;
  wire yshift_26__ap_start;
  wire yshift_26__ap_ready;
  wire yshift_26__ap_done;
  wire yshift_26__ap_idle;
  reg [1:0] yshift_26__state;
  reg [1:0] tapa_state;
  reg [0:0] countdown;
  wire ap_start__q0;
  wire ap_done__q0;
  assign Mmap2Stream_0___n__q0 = n;
  assign Mmap2Stream_0___rmem0__q0 = rmem0;
  assign Mmap2Stream_0__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_0__is_done__q0 = (Mmap2Stream_0__state == 2'b10);
  assign Mmap2Stream_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_0__state <= 2'b00;
    end else begin
      if(Mmap2Stream_0__state == 2'b00) begin
        if(Mmap2Stream_0__ap_start_global__q0) begin
          Mmap2Stream_0__state <= 2'b01;
        end 
      end 
      if(Mmap2Stream_0__state == 2'b01) begin
        if(Mmap2Stream_0__ap_ready) begin
          if(Mmap2Stream_0__ap_done) begin
            Mmap2Stream_0__state <= 2'b10;
          end else begin
            Mmap2Stream_0__state <= 2'b11;
          end
        end 
      end 
      if(Mmap2Stream_0__state == 2'b11) begin
        if(Mmap2Stream_0__ap_done) begin
          Mmap2Stream_0__state <= 2'b10;
        end 
      end 
      if(Mmap2Stream_0__state == 2'b10) begin
        if(Mmap2Stream_0__ap_done_global__q0) begin
          Mmap2Stream_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign Mmap2Stream_0__ap_start = (Mmap2Stream_0__state == 2'b01);
  assign Mmap2Stream_1___n__q0 = n;
  assign Mmap2Stream_1___rmem1__q0 = rmem1;
  assign Mmap2Stream_1__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_1__is_done__q0 = (Mmap2Stream_1__state == 2'b10);
  assign Mmap2Stream_1__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_1__state <= 2'b00;
    end else begin
      if(Mmap2Stream_1__state == 2'b00) begin
        if(Mmap2Stream_1__ap_start_global__q0) begin
          Mmap2Stream_1__state <= 2'b01;
        end 
      end 
      if(Mmap2Stream_1__state == 2'b01) begin
        if(Mmap2Stream_1__ap_ready) begin
          if(Mmap2Stream_1__ap_done) begin
            Mmap2Stream_1__state <= 2'b10;
          end else begin
            Mmap2Stream_1__state <= 2'b11;
          end
        end 
      end 
      if(Mmap2Stream_1__state == 2'b11) begin
        if(Mmap2Stream_1__ap_done) begin
          Mmap2Stream_1__state <= 2'b10;
        end 
      end 
      if(Mmap2Stream_1__state == 2'b10) begin
        if(Mmap2Stream_1__ap_done_global__q0) begin
          Mmap2Stream_1__state <= 2'b00;
        end 
      end 
    end
  end

  assign Mmap2Stream_1__ap_start = (Mmap2Stream_1__state == 2'b01);
  assign Mmap2Stream_2___n__q0 = n;
  assign Mmap2Stream_2___rmem2__q0 = rmem2;
  assign Mmap2Stream_2__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_2__is_done__q0 = (Mmap2Stream_2__state == 2'b10);
  assign Mmap2Stream_2__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_2__state <= 2'b00;
    end else begin
      if(Mmap2Stream_2__state == 2'b00) begin
        if(Mmap2Stream_2__ap_start_global__q0) begin
          Mmap2Stream_2__state <= 2'b01;
        end 
      end 
      if(Mmap2Stream_2__state == 2'b01) begin
        if(Mmap2Stream_2__ap_ready) begin
          if(Mmap2Stream_2__ap_done) begin
            Mmap2Stream_2__state <= 2'b10;
          end else begin
            Mmap2Stream_2__state <= 2'b11;
          end
        end 
      end 
      if(Mmap2Stream_2__state == 2'b11) begin
        if(Mmap2Stream_2__ap_done) begin
          Mmap2Stream_2__state <= 2'b10;
        end 
      end 
      if(Mmap2Stream_2__state == 2'b10) begin
        if(Mmap2Stream_2__ap_done_global__q0) begin
          Mmap2Stream_2__state <= 2'b00;
        end 
      end 
    end
  end

  assign Mmap2Stream_2__ap_start = (Mmap2Stream_2__state == 2'b01);
  assign Mmap2Stream_3___n__q0 = n;
  assign Mmap2Stream_3___rmem3__q0 = rmem3;
  assign Mmap2Stream_3__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_3__is_done__q0 = (Mmap2Stream_3__state == 2'b10);
  assign Mmap2Stream_3__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_3__state <= 2'b00;
    end else begin
      if(Mmap2Stream_3__state == 2'b00) begin
        if(Mmap2Stream_3__ap_start_global__q0) begin
          Mmap2Stream_3__state <= 2'b01;
        end 
      end 
      if(Mmap2Stream_3__state == 2'b01) begin
        if(Mmap2Stream_3__ap_ready) begin
          if(Mmap2Stream_3__ap_done) begin
            Mmap2Stream_3__state <= 2'b10;
          end else begin
            Mmap2Stream_3__state <= 2'b11;
          end
        end 
      end 
      if(Mmap2Stream_3__state == 2'b11) begin
        if(Mmap2Stream_3__ap_done) begin
          Mmap2Stream_3__state <= 2'b10;
        end 
      end 
      if(Mmap2Stream_3__state == 2'b10) begin
        if(Mmap2Stream_3__ap_done_global__q0) begin
          Mmap2Stream_3__state <= 2'b00;
        end 
      end 
    end
  end

  assign Mmap2Stream_3__ap_start = (Mmap2Stream_3__state == 2'b01);
  assign Mmap2Stream_4___n__q0 = n;
  assign Mmap2Stream_4___rmem4__q0 = rmem4;
  assign Mmap2Stream_4__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_4__is_done__q0 = (Mmap2Stream_4__state == 2'b10);
  assign Mmap2Stream_4__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_4__state <= 2'b00;
    end else begin
      if(Mmap2Stream_4__state == 2'b00) begin
        if(Mmap2Stream_4__ap_start_global__q0) begin
          Mmap2Stream_4__state <= 2'b01;
        end 
      end 
      if(Mmap2Stream_4__state == 2'b01) begin
        if(Mmap2Stream_4__ap_ready) begin
          if(Mmap2Stream_4__ap_done) begin
            Mmap2Stream_4__state <= 2'b10;
          end else begin
            Mmap2Stream_4__state <= 2'b11;
          end
        end 
      end 
      if(Mmap2Stream_4__state == 2'b11) begin
        if(Mmap2Stream_4__ap_done) begin
          Mmap2Stream_4__state <= 2'b10;
        end 
      end 
      if(Mmap2Stream_4__state == 2'b10) begin
        if(Mmap2Stream_4__ap_done_global__q0) begin
          Mmap2Stream_4__state <= 2'b00;
        end 
      end 
    end
  end

  assign Mmap2Stream_4__ap_start = (Mmap2Stream_4__state == 2'b01);
  assign Mmap2Stream_5___n__q0 = n;
  assign Mmap2Stream_5___rmem5__q0 = rmem5;
  assign Mmap2Stream_5__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_5__is_done__q0 = (Mmap2Stream_5__state == 2'b10);
  assign Mmap2Stream_5__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_5__state <= 2'b00;
    end else begin
      if(Mmap2Stream_5__state == 2'b00) begin
        if(Mmap2Stream_5__ap_start_global__q0) begin
          Mmap2Stream_5__state <= 2'b01;
        end 
      end 
      if(Mmap2Stream_5__state == 2'b01) begin
        if(Mmap2Stream_5__ap_ready) begin
          if(Mmap2Stream_5__ap_done) begin
            Mmap2Stream_5__state <= 2'b10;
          end else begin
            Mmap2Stream_5__state <= 2'b11;
          end
        end 
      end 
      if(Mmap2Stream_5__state == 2'b11) begin
        if(Mmap2Stream_5__ap_done) begin
          Mmap2Stream_5__state <= 2'b10;
        end 
      end 
      if(Mmap2Stream_5__state == 2'b10) begin
        if(Mmap2Stream_5__ap_done_global__q0) begin
          Mmap2Stream_5__state <= 2'b00;
        end 
      end 
    end
  end

  assign Mmap2Stream_5__ap_start = (Mmap2Stream_5__state == 2'b01);
  assign Mmap2Stream_6___n__q0 = n;
  assign Mmap2Stream_6___rmem6__q0 = rmem6;
  assign Mmap2Stream_6__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_6__is_done__q0 = (Mmap2Stream_6__state == 2'b10);
  assign Mmap2Stream_6__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_6__state <= 2'b00;
    end else begin
      if(Mmap2Stream_6__state == 2'b00) begin
        if(Mmap2Stream_6__ap_start_global__q0) begin
          Mmap2Stream_6__state <= 2'b01;
        end 
      end 
      if(Mmap2Stream_6__state == 2'b01) begin
        if(Mmap2Stream_6__ap_ready) begin
          if(Mmap2Stream_6__ap_done) begin
            Mmap2Stream_6__state <= 2'b10;
          end else begin
            Mmap2Stream_6__state <= 2'b11;
          end
        end 
      end 
      if(Mmap2Stream_6__state == 2'b11) begin
        if(Mmap2Stream_6__ap_done) begin
          Mmap2Stream_6__state <= 2'b10;
        end 
      end 
      if(Mmap2Stream_6__state == 2'b10) begin
        if(Mmap2Stream_6__ap_done_global__q0) begin
          Mmap2Stream_6__state <= 2'b00;
        end 
      end 
    end
  end

  assign Mmap2Stream_6__ap_start = (Mmap2Stream_6__state == 2'b01);
  assign Mmap2Stream_7___n__q0 = n;
  assign Mmap2Stream_7___rmem7__q0 = rmem7;
  assign Mmap2Stream_7__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_7__is_done__q0 = (Mmap2Stream_7__state == 2'b10);
  assign Mmap2Stream_7__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_7__state <= 2'b00;
    end else begin
      if(Mmap2Stream_7__state == 2'b00) begin
        if(Mmap2Stream_7__ap_start_global__q0) begin
          Mmap2Stream_7__state <= 2'b01;
        end 
      end 
      if(Mmap2Stream_7__state == 2'b01) begin
        if(Mmap2Stream_7__ap_ready) begin
          if(Mmap2Stream_7__ap_done) begin
            Mmap2Stream_7__state <= 2'b10;
          end else begin
            Mmap2Stream_7__state <= 2'b11;
          end
        end 
      end 
      if(Mmap2Stream_7__state == 2'b11) begin
        if(Mmap2Stream_7__ap_done) begin
          Mmap2Stream_7__state <= 2'b10;
        end 
      end 
      if(Mmap2Stream_7__state == 2'b10) begin
        if(Mmap2Stream_7__ap_done_global__q0) begin
          Mmap2Stream_7__state <= 2'b00;
        end 
      end 
    end
  end

  assign Mmap2Stream_7__ap_start = (Mmap2Stream_7__state == 2'b01);
  assign Mmap2Stream_8___n__q0 = n;
  assign Mmap2Stream_8___rmem8__q0 = rmem8;
  assign Mmap2Stream_8__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_8__is_done__q0 = (Mmap2Stream_8__state == 2'b10);
  assign Mmap2Stream_8__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_8__state <= 2'b00;
    end else begin
      if(Mmap2Stream_8__state == 2'b00) begin
        if(Mmap2Stream_8__ap_start_global__q0) begin
          Mmap2Stream_8__state <= 2'b01;
        end 
      end 
      if(Mmap2Stream_8__state == 2'b01) begin
        if(Mmap2Stream_8__ap_ready) begin
          if(Mmap2Stream_8__ap_done) begin
            Mmap2Stream_8__state <= 2'b10;
          end else begin
            Mmap2Stream_8__state <= 2'b11;
          end
        end 
      end 
      if(Mmap2Stream_8__state == 2'b11) begin
        if(Mmap2Stream_8__ap_done) begin
          Mmap2Stream_8__state <= 2'b10;
        end 
      end 
      if(Mmap2Stream_8__state == 2'b10) begin
        if(Mmap2Stream_8__ap_done_global__q0) begin
          Mmap2Stream_8__state <= 2'b00;
        end 
      end 
    end
  end

  assign Mmap2Stream_8__ap_start = (Mmap2Stream_8__state == 2'b01);
  assign Mmap2Stream_9___n__q0 = n;
  assign Mmap2Stream_9___rmem9__q0 = rmem9;
  assign Mmap2Stream_9__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_9__is_done__q0 = (Mmap2Stream_9__state == 2'b10);
  assign Mmap2Stream_9__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_9__state <= 2'b00;
    end else begin
      if(Mmap2Stream_9__state == 2'b00) begin
        if(Mmap2Stream_9__ap_start_global__q0) begin
          Mmap2Stream_9__state <= 2'b01;
        end 
      end 
      if(Mmap2Stream_9__state == 2'b01) begin
        if(Mmap2Stream_9__ap_ready) begin
          if(Mmap2Stream_9__ap_done) begin
            Mmap2Stream_9__state <= 2'b10;
          end else begin
            Mmap2Stream_9__state <= 2'b11;
          end
        end 
      end 
      if(Mmap2Stream_9__state == 2'b11) begin
        if(Mmap2Stream_9__ap_done) begin
          Mmap2Stream_9__state <= 2'b10;
        end 
      end 
      if(Mmap2Stream_9__state == 2'b10) begin
        if(Mmap2Stream_9__ap_done_global__q0) begin
          Mmap2Stream_9__state <= 2'b00;
        end 
      end 
    end
  end

  assign Mmap2Stream_9__ap_start = (Mmap2Stream_9__state == 2'b01);
  assign Mmap2Stream_10___n__q0 = n;
  assign Mmap2Stream_10___rmem10__q0 = rmem10;
  assign Mmap2Stream_10__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_10__is_done__q0 = (Mmap2Stream_10__state == 2'b10);
  assign Mmap2Stream_10__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_10__state <= 2'b00;
    end else begin
      if(Mmap2Stream_10__state == 2'b00) begin
        if(Mmap2Stream_10__ap_start_global__q0) begin
          Mmap2Stream_10__state <= 2'b01;
        end 
      end 
      if(Mmap2Stream_10__state == 2'b01) begin
        if(Mmap2Stream_10__ap_ready) begin
          if(Mmap2Stream_10__ap_done) begin
            Mmap2Stream_10__state <= 2'b10;
          end else begin
            Mmap2Stream_10__state <= 2'b11;
          end
        end 
      end 
      if(Mmap2Stream_10__state == 2'b11) begin
        if(Mmap2Stream_10__ap_done) begin
          Mmap2Stream_10__state <= 2'b10;
        end 
      end 
      if(Mmap2Stream_10__state == 2'b10) begin
        if(Mmap2Stream_10__ap_done_global__q0) begin
          Mmap2Stream_10__state <= 2'b00;
        end 
      end 
    end
  end

  assign Mmap2Stream_10__ap_start = (Mmap2Stream_10__state == 2'b01);
  assign Mmap2Stream_11___n__q0 = n;
  assign Mmap2Stream_11___rmem11__q0 = rmem11;
  assign Mmap2Stream_11__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_11__is_done__q0 = (Mmap2Stream_11__state == 2'b10);
  assign Mmap2Stream_11__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_11__state <= 2'b00;
    end else begin
      if(Mmap2Stream_11__state == 2'b00) begin
        if(Mmap2Stream_11__ap_start_global__q0) begin
          Mmap2Stream_11__state <= 2'b01;
        end 
      end 
      if(Mmap2Stream_11__state == 2'b01) begin
        if(Mmap2Stream_11__ap_ready) begin
          if(Mmap2Stream_11__ap_done) begin
            Mmap2Stream_11__state <= 2'b10;
          end else begin
            Mmap2Stream_11__state <= 2'b11;
          end
        end 
      end 
      if(Mmap2Stream_11__state == 2'b11) begin
        if(Mmap2Stream_11__ap_done) begin
          Mmap2Stream_11__state <= 2'b10;
        end 
      end 
      if(Mmap2Stream_11__state == 2'b10) begin
        if(Mmap2Stream_11__ap_done_global__q0) begin
          Mmap2Stream_11__state <= 2'b00;
        end 
      end 
    end
  end

  assign Mmap2Stream_11__ap_start = (Mmap2Stream_11__state == 2'b01);
  assign Mmap2Stream_12___n__q0 = n;
  assign Mmap2Stream_12___rmem12__q0 = rmem12;
  assign Mmap2Stream_12__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_12__is_done__q0 = (Mmap2Stream_12__state == 2'b10);
  assign Mmap2Stream_12__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_12__state <= 2'b00;
    end else begin
      if(Mmap2Stream_12__state == 2'b00) begin
        if(Mmap2Stream_12__ap_start_global__q0) begin
          Mmap2Stream_12__state <= 2'b01;
        end 
      end 
      if(Mmap2Stream_12__state == 2'b01) begin
        if(Mmap2Stream_12__ap_ready) begin
          if(Mmap2Stream_12__ap_done) begin
            Mmap2Stream_12__state <= 2'b10;
          end else begin
            Mmap2Stream_12__state <= 2'b11;
          end
        end 
      end 
      if(Mmap2Stream_12__state == 2'b11) begin
        if(Mmap2Stream_12__ap_done) begin
          Mmap2Stream_12__state <= 2'b10;
        end 
      end 
      if(Mmap2Stream_12__state == 2'b10) begin
        if(Mmap2Stream_12__ap_done_global__q0) begin
          Mmap2Stream_12__state <= 2'b00;
        end 
      end 
    end
  end

  assign Mmap2Stream_12__ap_start = (Mmap2Stream_12__state == 2'b01);
  assign Mmap2Stream_13___n__q0 = n;
  assign Mmap2Stream_13___rmem13__q0 = rmem13;
  assign Mmap2Stream_13__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_13__is_done__q0 = (Mmap2Stream_13__state == 2'b10);
  assign Mmap2Stream_13__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_13__state <= 2'b00;
    end else begin
      if(Mmap2Stream_13__state == 2'b00) begin
        if(Mmap2Stream_13__ap_start_global__q0) begin
          Mmap2Stream_13__state <= 2'b01;
        end 
      end 
      if(Mmap2Stream_13__state == 2'b01) begin
        if(Mmap2Stream_13__ap_ready) begin
          if(Mmap2Stream_13__ap_done) begin
            Mmap2Stream_13__state <= 2'b10;
          end else begin
            Mmap2Stream_13__state <= 2'b11;
          end
        end 
      end 
      if(Mmap2Stream_13__state == 2'b11) begin
        if(Mmap2Stream_13__ap_done) begin
          Mmap2Stream_13__state <= 2'b10;
        end 
      end 
      if(Mmap2Stream_13__state == 2'b10) begin
        if(Mmap2Stream_13__ap_done_global__q0) begin
          Mmap2Stream_13__state <= 2'b00;
        end 
      end 
    end
  end

  assign Mmap2Stream_13__ap_start = (Mmap2Stream_13__state == 2'b01);
  assign Mmap2Stream_14___n__q0 = n;
  assign Mmap2Stream_14___rmem14__q0 = rmem14;
  assign Mmap2Stream_14__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_14__is_done__q0 = (Mmap2Stream_14__state == 2'b10);
  assign Mmap2Stream_14__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_14__state <= 2'b00;
    end else begin
      if(Mmap2Stream_14__state == 2'b00) begin
        if(Mmap2Stream_14__ap_start_global__q0) begin
          Mmap2Stream_14__state <= 2'b01;
        end 
      end 
      if(Mmap2Stream_14__state == 2'b01) begin
        if(Mmap2Stream_14__ap_ready) begin
          if(Mmap2Stream_14__ap_done) begin
            Mmap2Stream_14__state <= 2'b10;
          end else begin
            Mmap2Stream_14__state <= 2'b11;
          end
        end 
      end 
      if(Mmap2Stream_14__state == 2'b11) begin
        if(Mmap2Stream_14__ap_done) begin
          Mmap2Stream_14__state <= 2'b10;
        end 
      end 
      if(Mmap2Stream_14__state == 2'b10) begin
        if(Mmap2Stream_14__ap_done_global__q0) begin
          Mmap2Stream_14__state <= 2'b00;
        end 
      end 
    end
  end

  assign Mmap2Stream_14__ap_start = (Mmap2Stream_14__state == 2'b01);
  assign Mmap2Stream_15___n__q0 = n;
  assign Mmap2Stream_15___rmem15__q0 = rmem15;
  assign Mmap2Stream_15__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_15__is_done__q0 = (Mmap2Stream_15__state == 2'b10);
  assign Mmap2Stream_15__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_15__state <= 2'b00;
    end else begin
      if(Mmap2Stream_15__state == 2'b00) begin
        if(Mmap2Stream_15__ap_start_global__q0) begin
          Mmap2Stream_15__state <= 2'b01;
        end 
      end 
      if(Mmap2Stream_15__state == 2'b01) begin
        if(Mmap2Stream_15__ap_ready) begin
          if(Mmap2Stream_15__ap_done) begin
            Mmap2Stream_15__state <= 2'b10;
          end else begin
            Mmap2Stream_15__state <= 2'b11;
          end
        end 
      end 
      if(Mmap2Stream_15__state == 2'b11) begin
        if(Mmap2Stream_15__ap_done) begin
          Mmap2Stream_15__state <= 2'b10;
        end 
      end 
      if(Mmap2Stream_15__state == 2'b10) begin
        if(Mmap2Stream_15__ap_done_global__q0) begin
          Mmap2Stream_15__state <= 2'b00;
        end 
      end 
    end
  end

  assign Mmap2Stream_15__ap_start = (Mmap2Stream_15__state == 2'b01);
  assign Mmap2Stream_16___n__q0 = n;
  assign Mmap2Stream_16___rmem16__q0 = rmem16;
  assign Mmap2Stream_16__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_16__is_done__q0 = (Mmap2Stream_16__state == 2'b10);
  assign Mmap2Stream_16__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_16__state <= 2'b00;
    end else begin
      if(Mmap2Stream_16__state == 2'b00) begin
        if(Mmap2Stream_16__ap_start_global__q0) begin
          Mmap2Stream_16__state <= 2'b01;
        end 
      end 
      if(Mmap2Stream_16__state == 2'b01) begin
        if(Mmap2Stream_16__ap_ready) begin
          if(Mmap2Stream_16__ap_done) begin
            Mmap2Stream_16__state <= 2'b10;
          end else begin
            Mmap2Stream_16__state <= 2'b11;
          end
        end 
      end 
      if(Mmap2Stream_16__state == 2'b11) begin
        if(Mmap2Stream_16__ap_done) begin
          Mmap2Stream_16__state <= 2'b10;
        end 
      end 
      if(Mmap2Stream_16__state == 2'b10) begin
        if(Mmap2Stream_16__ap_done_global__q0) begin
          Mmap2Stream_16__state <= 2'b00;
        end 
      end 
    end
  end

  assign Mmap2Stream_16__ap_start = (Mmap2Stream_16__state == 2'b01);
  assign Mmap2Stream_17___n__q0 = n;
  assign Mmap2Stream_17___rmem17__q0 = rmem17;
  assign Mmap2Stream_17__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_17__is_done__q0 = (Mmap2Stream_17__state == 2'b10);
  assign Mmap2Stream_17__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_17__state <= 2'b00;
    end else begin
      if(Mmap2Stream_17__state == 2'b00) begin
        if(Mmap2Stream_17__ap_start_global__q0) begin
          Mmap2Stream_17__state <= 2'b01;
        end 
      end 
      if(Mmap2Stream_17__state == 2'b01) begin
        if(Mmap2Stream_17__ap_ready) begin
          if(Mmap2Stream_17__ap_done) begin
            Mmap2Stream_17__state <= 2'b10;
          end else begin
            Mmap2Stream_17__state <= 2'b11;
          end
        end 
      end 
      if(Mmap2Stream_17__state == 2'b11) begin
        if(Mmap2Stream_17__ap_done) begin
          Mmap2Stream_17__state <= 2'b10;
        end 
      end 
      if(Mmap2Stream_17__state == 2'b10) begin
        if(Mmap2Stream_17__ap_done_global__q0) begin
          Mmap2Stream_17__state <= 2'b00;
        end 
      end 
    end
  end

  assign Mmap2Stream_17__ap_start = (Mmap2Stream_17__state == 2'b01);
  assign Mmap2Stream_18___n__q0 = n;
  assign Mmap2Stream_18___rmem18__q0 = rmem18;
  assign Mmap2Stream_18__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_18__is_done__q0 = (Mmap2Stream_18__state == 2'b10);
  assign Mmap2Stream_18__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_18__state <= 2'b00;
    end else begin
      if(Mmap2Stream_18__state == 2'b00) begin
        if(Mmap2Stream_18__ap_start_global__q0) begin
          Mmap2Stream_18__state <= 2'b01;
        end 
      end 
      if(Mmap2Stream_18__state == 2'b01) begin
        if(Mmap2Stream_18__ap_ready) begin
          if(Mmap2Stream_18__ap_done) begin
            Mmap2Stream_18__state <= 2'b10;
          end else begin
            Mmap2Stream_18__state <= 2'b11;
          end
        end 
      end 
      if(Mmap2Stream_18__state == 2'b11) begin
        if(Mmap2Stream_18__ap_done) begin
          Mmap2Stream_18__state <= 2'b10;
        end 
      end 
      if(Mmap2Stream_18__state == 2'b10) begin
        if(Mmap2Stream_18__ap_done_global__q0) begin
          Mmap2Stream_18__state <= 2'b00;
        end 
      end 
    end
  end

  assign Mmap2Stream_18__ap_start = (Mmap2Stream_18__state == 2'b01);
  assign Mmap2Stream_19___n__q0 = n;
  assign Mmap2Stream_19___rmem19__q0 = rmem19;
  assign Mmap2Stream_19__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_19__is_done__q0 = (Mmap2Stream_19__state == 2'b10);
  assign Mmap2Stream_19__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_19__state <= 2'b00;
    end else begin
      if(Mmap2Stream_19__state == 2'b00) begin
        if(Mmap2Stream_19__ap_start_global__q0) begin
          Mmap2Stream_19__state <= 2'b01;
        end 
      end 
      if(Mmap2Stream_19__state == 2'b01) begin
        if(Mmap2Stream_19__ap_ready) begin
          if(Mmap2Stream_19__ap_done) begin
            Mmap2Stream_19__state <= 2'b10;
          end else begin
            Mmap2Stream_19__state <= 2'b11;
          end
        end 
      end 
      if(Mmap2Stream_19__state == 2'b11) begin
        if(Mmap2Stream_19__ap_done) begin
          Mmap2Stream_19__state <= 2'b10;
        end 
      end 
      if(Mmap2Stream_19__state == 2'b10) begin
        if(Mmap2Stream_19__ap_done_global__q0) begin
          Mmap2Stream_19__state <= 2'b00;
        end 
      end 
    end
  end

  assign Mmap2Stream_19__ap_start = (Mmap2Stream_19__state == 2'b01);
  assign Mmap2Stream_20___n__q0 = n;
  assign Mmap2Stream_20___rmem20__q0 = rmem20;
  assign Mmap2Stream_20__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_20__is_done__q0 = (Mmap2Stream_20__state == 2'b10);
  assign Mmap2Stream_20__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_20__state <= 2'b00;
    end else begin
      if(Mmap2Stream_20__state == 2'b00) begin
        if(Mmap2Stream_20__ap_start_global__q0) begin
          Mmap2Stream_20__state <= 2'b01;
        end 
      end 
      if(Mmap2Stream_20__state == 2'b01) begin
        if(Mmap2Stream_20__ap_ready) begin
          if(Mmap2Stream_20__ap_done) begin
            Mmap2Stream_20__state <= 2'b10;
          end else begin
            Mmap2Stream_20__state <= 2'b11;
          end
        end 
      end 
      if(Mmap2Stream_20__state == 2'b11) begin
        if(Mmap2Stream_20__ap_done) begin
          Mmap2Stream_20__state <= 2'b10;
        end 
      end 
      if(Mmap2Stream_20__state == 2'b10) begin
        if(Mmap2Stream_20__ap_done_global__q0) begin
          Mmap2Stream_20__state <= 2'b00;
        end 
      end 
    end
  end

  assign Mmap2Stream_20__ap_start = (Mmap2Stream_20__state == 2'b01);
  assign Mmap2Stream_21___n__q0 = n;
  assign Mmap2Stream_21___rmem21__q0 = rmem21;
  assign Mmap2Stream_21__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_21__is_done__q0 = (Mmap2Stream_21__state == 2'b10);
  assign Mmap2Stream_21__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_21__state <= 2'b00;
    end else begin
      if(Mmap2Stream_21__state == 2'b00) begin
        if(Mmap2Stream_21__ap_start_global__q0) begin
          Mmap2Stream_21__state <= 2'b01;
        end 
      end 
      if(Mmap2Stream_21__state == 2'b01) begin
        if(Mmap2Stream_21__ap_ready) begin
          if(Mmap2Stream_21__ap_done) begin
            Mmap2Stream_21__state <= 2'b10;
          end else begin
            Mmap2Stream_21__state <= 2'b11;
          end
        end 
      end 
      if(Mmap2Stream_21__state == 2'b11) begin
        if(Mmap2Stream_21__ap_done) begin
          Mmap2Stream_21__state <= 2'b10;
        end 
      end 
      if(Mmap2Stream_21__state == 2'b10) begin
        if(Mmap2Stream_21__ap_done_global__q0) begin
          Mmap2Stream_21__state <= 2'b00;
        end 
      end 
    end
  end

  assign Mmap2Stream_21__ap_start = (Mmap2Stream_21__state == 2'b01);
  assign Mmap2Stream_22___n__q0 = n;
  assign Mmap2Stream_22___rmem22__q0 = rmem22;
  assign Mmap2Stream_22__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_22__is_done__q0 = (Mmap2Stream_22__state == 2'b10);
  assign Mmap2Stream_22__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_22__state <= 2'b00;
    end else begin
      if(Mmap2Stream_22__state == 2'b00) begin
        if(Mmap2Stream_22__ap_start_global__q0) begin
          Mmap2Stream_22__state <= 2'b01;
        end 
      end 
      if(Mmap2Stream_22__state == 2'b01) begin
        if(Mmap2Stream_22__ap_ready) begin
          if(Mmap2Stream_22__ap_done) begin
            Mmap2Stream_22__state <= 2'b10;
          end else begin
            Mmap2Stream_22__state <= 2'b11;
          end
        end 
      end 
      if(Mmap2Stream_22__state == 2'b11) begin
        if(Mmap2Stream_22__ap_done) begin
          Mmap2Stream_22__state <= 2'b10;
        end 
      end 
      if(Mmap2Stream_22__state == 2'b10) begin
        if(Mmap2Stream_22__ap_done_global__q0) begin
          Mmap2Stream_22__state <= 2'b00;
        end 
      end 
    end
  end

  assign Mmap2Stream_22__ap_start = (Mmap2Stream_22__state == 2'b01);
  assign Mmap2Stream_23___n__q0 = n;
  assign Mmap2Stream_23___rmem23__q0 = rmem23;
  assign Mmap2Stream_23__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_23__is_done__q0 = (Mmap2Stream_23__state == 2'b10);
  assign Mmap2Stream_23__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_23__state <= 2'b00;
    end else begin
      if(Mmap2Stream_23__state == 2'b00) begin
        if(Mmap2Stream_23__ap_start_global__q0) begin
          Mmap2Stream_23__state <= 2'b01;
        end 
      end 
      if(Mmap2Stream_23__state == 2'b01) begin
        if(Mmap2Stream_23__ap_ready) begin
          if(Mmap2Stream_23__ap_done) begin
            Mmap2Stream_23__state <= 2'b10;
          end else begin
            Mmap2Stream_23__state <= 2'b11;
          end
        end 
      end 
      if(Mmap2Stream_23__state == 2'b11) begin
        if(Mmap2Stream_23__ap_done) begin
          Mmap2Stream_23__state <= 2'b10;
        end 
      end 
      if(Mmap2Stream_23__state == 2'b10) begin
        if(Mmap2Stream_23__ap_done_global__q0) begin
          Mmap2Stream_23__state <= 2'b00;
        end 
      end 
    end
  end

  assign Mmap2Stream_23__ap_start = (Mmap2Stream_23__state == 2'b01);
  assign Mmap2Stream_24___n__q0 = n;
  assign Mmap2Stream_24___rmem24__q0 = rmem24;
  assign Mmap2Stream_24__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_24__is_done__q0 = (Mmap2Stream_24__state == 2'b10);
  assign Mmap2Stream_24__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_24__state <= 2'b00;
    end else begin
      if(Mmap2Stream_24__state == 2'b00) begin
        if(Mmap2Stream_24__ap_start_global__q0) begin
          Mmap2Stream_24__state <= 2'b01;
        end 
      end 
      if(Mmap2Stream_24__state == 2'b01) begin
        if(Mmap2Stream_24__ap_ready) begin
          if(Mmap2Stream_24__ap_done) begin
            Mmap2Stream_24__state <= 2'b10;
          end else begin
            Mmap2Stream_24__state <= 2'b11;
          end
        end 
      end 
      if(Mmap2Stream_24__state == 2'b11) begin
        if(Mmap2Stream_24__ap_done) begin
          Mmap2Stream_24__state <= 2'b10;
        end 
      end 
      if(Mmap2Stream_24__state == 2'b10) begin
        if(Mmap2Stream_24__ap_done_global__q0) begin
          Mmap2Stream_24__state <= 2'b00;
        end 
      end 
    end
  end

  assign Mmap2Stream_24__ap_start = (Mmap2Stream_24__state == 2'b01);
  assign Mmap2Stream_25___n__q0 = n;
  assign Mmap2Stream_25___rmem25__q0 = rmem25;
  assign Mmap2Stream_25__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_25__is_done__q0 = (Mmap2Stream_25__state == 2'b10);
  assign Mmap2Stream_25__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_25__state <= 2'b00;
    end else begin
      if(Mmap2Stream_25__state == 2'b00) begin
        if(Mmap2Stream_25__ap_start_global__q0) begin
          Mmap2Stream_25__state <= 2'b01;
        end 
      end 
      if(Mmap2Stream_25__state == 2'b01) begin
        if(Mmap2Stream_25__ap_ready) begin
          if(Mmap2Stream_25__ap_done) begin
            Mmap2Stream_25__state <= 2'b10;
          end else begin
            Mmap2Stream_25__state <= 2'b11;
          end
        end 
      end 
      if(Mmap2Stream_25__state == 2'b11) begin
        if(Mmap2Stream_25__ap_done) begin
          Mmap2Stream_25__state <= 2'b10;
        end 
      end 
      if(Mmap2Stream_25__state == 2'b10) begin
        if(Mmap2Stream_25__ap_done_global__q0) begin
          Mmap2Stream_25__state <= 2'b00;
        end 
      end 
    end
  end

  assign Mmap2Stream_25__ap_start = (Mmap2Stream_25__state == 2'b01);
  assign Mmap2Stream_26___n__q0 = n;
  assign Mmap2Stream_26___rmem26__q0 = rmem26;
  assign Mmap2Stream_26__ap_start_global__q0 = ap_start__q0;
  assign Mmap2Stream_26__is_done__q0 = (Mmap2Stream_26__state == 2'b10);
  assign Mmap2Stream_26__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Mmap2Stream_26__state <= 2'b00;
    end else begin
      if(Mmap2Stream_26__state == 2'b00) begin
        if(Mmap2Stream_26__ap_start_global__q0) begin
          Mmap2Stream_26__state <= 2'b01;
        end 
      end 
      if(Mmap2Stream_26__state == 2'b01) begin
        if(Mmap2Stream_26__ap_ready) begin
          if(Mmap2Stream_26__ap_done) begin
            Mmap2Stream_26__state <= 2'b10;
          end else begin
            Mmap2Stream_26__state <= 2'b11;
          end
        end 
      end 
      if(Mmap2Stream_26__state == 2'b11) begin
        if(Mmap2Stream_26__ap_done) begin
          Mmap2Stream_26__state <= 2'b10;
        end 
      end 
      if(Mmap2Stream_26__state == 2'b10) begin
        if(Mmap2Stream_26__ap_done_global__q0) begin
          Mmap2Stream_26__state <= 2'b00;
        end 
      end 
    end
  end

  assign Mmap2Stream_26__ap_start = (Mmap2Stream_26__state == 2'b01);
  assign Stream2Mmap_0___n__q0 = n;
  assign Stream2Mmap_0___rmem0__q0 = rmem0;
  assign Stream2Mmap_0__ap_start_global__q0 = ap_start__q0;
  assign Stream2Mmap_0__is_done__q0 = (Stream2Mmap_0__state == 2'b10);
  assign Stream2Mmap_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Stream2Mmap_0__state <= 2'b00;
    end else begin
      if(Stream2Mmap_0__state == 2'b00) begin
        if(Stream2Mmap_0__ap_start_global__q0) begin
          Stream2Mmap_0__state <= 2'b01;
        end 
      end 
      if(Stream2Mmap_0__state == 2'b01) begin
        if(Stream2Mmap_0__ap_ready) begin
          if(Stream2Mmap_0__ap_done) begin
            Stream2Mmap_0__state <= 2'b10;
          end else begin
            Stream2Mmap_0__state <= 2'b11;
          end
        end 
      end 
      if(Stream2Mmap_0__state == 2'b11) begin
        if(Stream2Mmap_0__ap_done) begin
          Stream2Mmap_0__state <= 2'b10;
        end 
      end 
      if(Stream2Mmap_0__state == 2'b10) begin
        if(Stream2Mmap_0__ap_done_global__q0) begin
          Stream2Mmap_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign Stream2Mmap_0__ap_start = (Stream2Mmap_0__state == 2'b01);
  assign Stream2Mmap_1___n__q0 = n;
  assign Stream2Mmap_1___rmem1__q0 = rmem1;
  assign Stream2Mmap_1__ap_start_global__q0 = ap_start__q0;
  assign Stream2Mmap_1__is_done__q0 = (Stream2Mmap_1__state == 2'b10);
  assign Stream2Mmap_1__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Stream2Mmap_1__state <= 2'b00;
    end else begin
      if(Stream2Mmap_1__state == 2'b00) begin
        if(Stream2Mmap_1__ap_start_global__q0) begin
          Stream2Mmap_1__state <= 2'b01;
        end 
      end 
      if(Stream2Mmap_1__state == 2'b01) begin
        if(Stream2Mmap_1__ap_ready) begin
          if(Stream2Mmap_1__ap_done) begin
            Stream2Mmap_1__state <= 2'b10;
          end else begin
            Stream2Mmap_1__state <= 2'b11;
          end
        end 
      end 
      if(Stream2Mmap_1__state == 2'b11) begin
        if(Stream2Mmap_1__ap_done) begin
          Stream2Mmap_1__state <= 2'b10;
        end 
      end 
      if(Stream2Mmap_1__state == 2'b10) begin
        if(Stream2Mmap_1__ap_done_global__q0) begin
          Stream2Mmap_1__state <= 2'b00;
        end 
      end 
    end
  end

  assign Stream2Mmap_1__ap_start = (Stream2Mmap_1__state == 2'b01);
  assign Stream2Mmap_2___n__q0 = n;
  assign Stream2Mmap_2___rmem2__q0 = rmem2;
  assign Stream2Mmap_2__ap_start_global__q0 = ap_start__q0;
  assign Stream2Mmap_2__is_done__q0 = (Stream2Mmap_2__state == 2'b10);
  assign Stream2Mmap_2__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Stream2Mmap_2__state <= 2'b00;
    end else begin
      if(Stream2Mmap_2__state == 2'b00) begin
        if(Stream2Mmap_2__ap_start_global__q0) begin
          Stream2Mmap_2__state <= 2'b01;
        end 
      end 
      if(Stream2Mmap_2__state == 2'b01) begin
        if(Stream2Mmap_2__ap_ready) begin
          if(Stream2Mmap_2__ap_done) begin
            Stream2Mmap_2__state <= 2'b10;
          end else begin
            Stream2Mmap_2__state <= 2'b11;
          end
        end 
      end 
      if(Stream2Mmap_2__state == 2'b11) begin
        if(Stream2Mmap_2__ap_done) begin
          Stream2Mmap_2__state <= 2'b10;
        end 
      end 
      if(Stream2Mmap_2__state == 2'b10) begin
        if(Stream2Mmap_2__ap_done_global__q0) begin
          Stream2Mmap_2__state <= 2'b00;
        end 
      end 
    end
  end

  assign Stream2Mmap_2__ap_start = (Stream2Mmap_2__state == 2'b01);
  assign Stream2Mmap_3___n__q0 = n;
  assign Stream2Mmap_3___rmem3__q0 = rmem3;
  assign Stream2Mmap_3__ap_start_global__q0 = ap_start__q0;
  assign Stream2Mmap_3__is_done__q0 = (Stream2Mmap_3__state == 2'b10);
  assign Stream2Mmap_3__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Stream2Mmap_3__state <= 2'b00;
    end else begin
      if(Stream2Mmap_3__state == 2'b00) begin
        if(Stream2Mmap_3__ap_start_global__q0) begin
          Stream2Mmap_3__state <= 2'b01;
        end 
      end 
      if(Stream2Mmap_3__state == 2'b01) begin
        if(Stream2Mmap_3__ap_ready) begin
          if(Stream2Mmap_3__ap_done) begin
            Stream2Mmap_3__state <= 2'b10;
          end else begin
            Stream2Mmap_3__state <= 2'b11;
          end
        end 
      end 
      if(Stream2Mmap_3__state == 2'b11) begin
        if(Stream2Mmap_3__ap_done) begin
          Stream2Mmap_3__state <= 2'b10;
        end 
      end 
      if(Stream2Mmap_3__state == 2'b10) begin
        if(Stream2Mmap_3__ap_done_global__q0) begin
          Stream2Mmap_3__state <= 2'b00;
        end 
      end 
    end
  end

  assign Stream2Mmap_3__ap_start = (Stream2Mmap_3__state == 2'b01);
  assign Stream2Mmap_4___n__q0 = n;
  assign Stream2Mmap_4___rmem4__q0 = rmem4;
  assign Stream2Mmap_4__ap_start_global__q0 = ap_start__q0;
  assign Stream2Mmap_4__is_done__q0 = (Stream2Mmap_4__state == 2'b10);
  assign Stream2Mmap_4__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Stream2Mmap_4__state <= 2'b00;
    end else begin
      if(Stream2Mmap_4__state == 2'b00) begin
        if(Stream2Mmap_4__ap_start_global__q0) begin
          Stream2Mmap_4__state <= 2'b01;
        end 
      end 
      if(Stream2Mmap_4__state == 2'b01) begin
        if(Stream2Mmap_4__ap_ready) begin
          if(Stream2Mmap_4__ap_done) begin
            Stream2Mmap_4__state <= 2'b10;
          end else begin
            Stream2Mmap_4__state <= 2'b11;
          end
        end 
      end 
      if(Stream2Mmap_4__state == 2'b11) begin
        if(Stream2Mmap_4__ap_done) begin
          Stream2Mmap_4__state <= 2'b10;
        end 
      end 
      if(Stream2Mmap_4__state == 2'b10) begin
        if(Stream2Mmap_4__ap_done_global__q0) begin
          Stream2Mmap_4__state <= 2'b00;
        end 
      end 
    end
  end

  assign Stream2Mmap_4__ap_start = (Stream2Mmap_4__state == 2'b01);
  assign Stream2Mmap_5___n__q0 = n;
  assign Stream2Mmap_5___rmem5__q0 = rmem5;
  assign Stream2Mmap_5__ap_start_global__q0 = ap_start__q0;
  assign Stream2Mmap_5__is_done__q0 = (Stream2Mmap_5__state == 2'b10);
  assign Stream2Mmap_5__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Stream2Mmap_5__state <= 2'b00;
    end else begin
      if(Stream2Mmap_5__state == 2'b00) begin
        if(Stream2Mmap_5__ap_start_global__q0) begin
          Stream2Mmap_5__state <= 2'b01;
        end 
      end 
      if(Stream2Mmap_5__state == 2'b01) begin
        if(Stream2Mmap_5__ap_ready) begin
          if(Stream2Mmap_5__ap_done) begin
            Stream2Mmap_5__state <= 2'b10;
          end else begin
            Stream2Mmap_5__state <= 2'b11;
          end
        end 
      end 
      if(Stream2Mmap_5__state == 2'b11) begin
        if(Stream2Mmap_5__ap_done) begin
          Stream2Mmap_5__state <= 2'b10;
        end 
      end 
      if(Stream2Mmap_5__state == 2'b10) begin
        if(Stream2Mmap_5__ap_done_global__q0) begin
          Stream2Mmap_5__state <= 2'b00;
        end 
      end 
    end
  end

  assign Stream2Mmap_5__ap_start = (Stream2Mmap_5__state == 2'b01);
  assign Stream2Mmap_6___n__q0 = n;
  assign Stream2Mmap_6___rmem6__q0 = rmem6;
  assign Stream2Mmap_6__ap_start_global__q0 = ap_start__q0;
  assign Stream2Mmap_6__is_done__q0 = (Stream2Mmap_6__state == 2'b10);
  assign Stream2Mmap_6__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Stream2Mmap_6__state <= 2'b00;
    end else begin
      if(Stream2Mmap_6__state == 2'b00) begin
        if(Stream2Mmap_6__ap_start_global__q0) begin
          Stream2Mmap_6__state <= 2'b01;
        end 
      end 
      if(Stream2Mmap_6__state == 2'b01) begin
        if(Stream2Mmap_6__ap_ready) begin
          if(Stream2Mmap_6__ap_done) begin
            Stream2Mmap_6__state <= 2'b10;
          end else begin
            Stream2Mmap_6__state <= 2'b11;
          end
        end 
      end 
      if(Stream2Mmap_6__state == 2'b11) begin
        if(Stream2Mmap_6__ap_done) begin
          Stream2Mmap_6__state <= 2'b10;
        end 
      end 
      if(Stream2Mmap_6__state == 2'b10) begin
        if(Stream2Mmap_6__ap_done_global__q0) begin
          Stream2Mmap_6__state <= 2'b00;
        end 
      end 
    end
  end

  assign Stream2Mmap_6__ap_start = (Stream2Mmap_6__state == 2'b01);
  assign Stream2Mmap_7___n__q0 = n;
  assign Stream2Mmap_7___rmem7__q0 = rmem7;
  assign Stream2Mmap_7__ap_start_global__q0 = ap_start__q0;
  assign Stream2Mmap_7__is_done__q0 = (Stream2Mmap_7__state == 2'b10);
  assign Stream2Mmap_7__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Stream2Mmap_7__state <= 2'b00;
    end else begin
      if(Stream2Mmap_7__state == 2'b00) begin
        if(Stream2Mmap_7__ap_start_global__q0) begin
          Stream2Mmap_7__state <= 2'b01;
        end 
      end 
      if(Stream2Mmap_7__state == 2'b01) begin
        if(Stream2Mmap_7__ap_ready) begin
          if(Stream2Mmap_7__ap_done) begin
            Stream2Mmap_7__state <= 2'b10;
          end else begin
            Stream2Mmap_7__state <= 2'b11;
          end
        end 
      end 
      if(Stream2Mmap_7__state == 2'b11) begin
        if(Stream2Mmap_7__ap_done) begin
          Stream2Mmap_7__state <= 2'b10;
        end 
      end 
      if(Stream2Mmap_7__state == 2'b10) begin
        if(Stream2Mmap_7__ap_done_global__q0) begin
          Stream2Mmap_7__state <= 2'b00;
        end 
      end 
    end
  end

  assign Stream2Mmap_7__ap_start = (Stream2Mmap_7__state == 2'b01);
  assign Stream2Mmap_8___n__q0 = n;
  assign Stream2Mmap_8___rmem8__q0 = rmem8;
  assign Stream2Mmap_8__ap_start_global__q0 = ap_start__q0;
  assign Stream2Mmap_8__is_done__q0 = (Stream2Mmap_8__state == 2'b10);
  assign Stream2Mmap_8__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Stream2Mmap_8__state <= 2'b00;
    end else begin
      if(Stream2Mmap_8__state == 2'b00) begin
        if(Stream2Mmap_8__ap_start_global__q0) begin
          Stream2Mmap_8__state <= 2'b01;
        end 
      end 
      if(Stream2Mmap_8__state == 2'b01) begin
        if(Stream2Mmap_8__ap_ready) begin
          if(Stream2Mmap_8__ap_done) begin
            Stream2Mmap_8__state <= 2'b10;
          end else begin
            Stream2Mmap_8__state <= 2'b11;
          end
        end 
      end 
      if(Stream2Mmap_8__state == 2'b11) begin
        if(Stream2Mmap_8__ap_done) begin
          Stream2Mmap_8__state <= 2'b10;
        end 
      end 
      if(Stream2Mmap_8__state == 2'b10) begin
        if(Stream2Mmap_8__ap_done_global__q0) begin
          Stream2Mmap_8__state <= 2'b00;
        end 
      end 
    end
  end

  assign Stream2Mmap_8__ap_start = (Stream2Mmap_8__state == 2'b01);
  assign Stream2Mmap_9___n__q0 = n;
  assign Stream2Mmap_9___rmem9__q0 = rmem9;
  assign Stream2Mmap_9__ap_start_global__q0 = ap_start__q0;
  assign Stream2Mmap_9__is_done__q0 = (Stream2Mmap_9__state == 2'b10);
  assign Stream2Mmap_9__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Stream2Mmap_9__state <= 2'b00;
    end else begin
      if(Stream2Mmap_9__state == 2'b00) begin
        if(Stream2Mmap_9__ap_start_global__q0) begin
          Stream2Mmap_9__state <= 2'b01;
        end 
      end 
      if(Stream2Mmap_9__state == 2'b01) begin
        if(Stream2Mmap_9__ap_ready) begin
          if(Stream2Mmap_9__ap_done) begin
            Stream2Mmap_9__state <= 2'b10;
          end else begin
            Stream2Mmap_9__state <= 2'b11;
          end
        end 
      end 
      if(Stream2Mmap_9__state == 2'b11) begin
        if(Stream2Mmap_9__ap_done) begin
          Stream2Mmap_9__state <= 2'b10;
        end 
      end 
      if(Stream2Mmap_9__state == 2'b10) begin
        if(Stream2Mmap_9__ap_done_global__q0) begin
          Stream2Mmap_9__state <= 2'b00;
        end 
      end 
    end
  end

  assign Stream2Mmap_9__ap_start = (Stream2Mmap_9__state == 2'b01);
  assign Stream2Mmap_10___n__q0 = n;
  assign Stream2Mmap_10___rmem10__q0 = rmem10;
  assign Stream2Mmap_10__ap_start_global__q0 = ap_start__q0;
  assign Stream2Mmap_10__is_done__q0 = (Stream2Mmap_10__state == 2'b10);
  assign Stream2Mmap_10__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Stream2Mmap_10__state <= 2'b00;
    end else begin
      if(Stream2Mmap_10__state == 2'b00) begin
        if(Stream2Mmap_10__ap_start_global__q0) begin
          Stream2Mmap_10__state <= 2'b01;
        end 
      end 
      if(Stream2Mmap_10__state == 2'b01) begin
        if(Stream2Mmap_10__ap_ready) begin
          if(Stream2Mmap_10__ap_done) begin
            Stream2Mmap_10__state <= 2'b10;
          end else begin
            Stream2Mmap_10__state <= 2'b11;
          end
        end 
      end 
      if(Stream2Mmap_10__state == 2'b11) begin
        if(Stream2Mmap_10__ap_done) begin
          Stream2Mmap_10__state <= 2'b10;
        end 
      end 
      if(Stream2Mmap_10__state == 2'b10) begin
        if(Stream2Mmap_10__ap_done_global__q0) begin
          Stream2Mmap_10__state <= 2'b00;
        end 
      end 
    end
  end

  assign Stream2Mmap_10__ap_start = (Stream2Mmap_10__state == 2'b01);
  assign Stream2Mmap_11___n__q0 = n;
  assign Stream2Mmap_11___rmem11__q0 = rmem11;
  assign Stream2Mmap_11__ap_start_global__q0 = ap_start__q0;
  assign Stream2Mmap_11__is_done__q0 = (Stream2Mmap_11__state == 2'b10);
  assign Stream2Mmap_11__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Stream2Mmap_11__state <= 2'b00;
    end else begin
      if(Stream2Mmap_11__state == 2'b00) begin
        if(Stream2Mmap_11__ap_start_global__q0) begin
          Stream2Mmap_11__state <= 2'b01;
        end 
      end 
      if(Stream2Mmap_11__state == 2'b01) begin
        if(Stream2Mmap_11__ap_ready) begin
          if(Stream2Mmap_11__ap_done) begin
            Stream2Mmap_11__state <= 2'b10;
          end else begin
            Stream2Mmap_11__state <= 2'b11;
          end
        end 
      end 
      if(Stream2Mmap_11__state == 2'b11) begin
        if(Stream2Mmap_11__ap_done) begin
          Stream2Mmap_11__state <= 2'b10;
        end 
      end 
      if(Stream2Mmap_11__state == 2'b10) begin
        if(Stream2Mmap_11__ap_done_global__q0) begin
          Stream2Mmap_11__state <= 2'b00;
        end 
      end 
    end
  end

  assign Stream2Mmap_11__ap_start = (Stream2Mmap_11__state == 2'b01);
  assign Stream2Mmap_12___n__q0 = n;
  assign Stream2Mmap_12___rmem12__q0 = rmem12;
  assign Stream2Mmap_12__ap_start_global__q0 = ap_start__q0;
  assign Stream2Mmap_12__is_done__q0 = (Stream2Mmap_12__state == 2'b10);
  assign Stream2Mmap_12__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Stream2Mmap_12__state <= 2'b00;
    end else begin
      if(Stream2Mmap_12__state == 2'b00) begin
        if(Stream2Mmap_12__ap_start_global__q0) begin
          Stream2Mmap_12__state <= 2'b01;
        end 
      end 
      if(Stream2Mmap_12__state == 2'b01) begin
        if(Stream2Mmap_12__ap_ready) begin
          if(Stream2Mmap_12__ap_done) begin
            Stream2Mmap_12__state <= 2'b10;
          end else begin
            Stream2Mmap_12__state <= 2'b11;
          end
        end 
      end 
      if(Stream2Mmap_12__state == 2'b11) begin
        if(Stream2Mmap_12__ap_done) begin
          Stream2Mmap_12__state <= 2'b10;
        end 
      end 
      if(Stream2Mmap_12__state == 2'b10) begin
        if(Stream2Mmap_12__ap_done_global__q0) begin
          Stream2Mmap_12__state <= 2'b00;
        end 
      end 
    end
  end

  assign Stream2Mmap_12__ap_start = (Stream2Mmap_12__state == 2'b01);
  assign Stream2Mmap_13___n__q0 = n;
  assign Stream2Mmap_13___rmem13__q0 = rmem13;
  assign Stream2Mmap_13__ap_start_global__q0 = ap_start__q0;
  assign Stream2Mmap_13__is_done__q0 = (Stream2Mmap_13__state == 2'b10);
  assign Stream2Mmap_13__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Stream2Mmap_13__state <= 2'b00;
    end else begin
      if(Stream2Mmap_13__state == 2'b00) begin
        if(Stream2Mmap_13__ap_start_global__q0) begin
          Stream2Mmap_13__state <= 2'b01;
        end 
      end 
      if(Stream2Mmap_13__state == 2'b01) begin
        if(Stream2Mmap_13__ap_ready) begin
          if(Stream2Mmap_13__ap_done) begin
            Stream2Mmap_13__state <= 2'b10;
          end else begin
            Stream2Mmap_13__state <= 2'b11;
          end
        end 
      end 
      if(Stream2Mmap_13__state == 2'b11) begin
        if(Stream2Mmap_13__ap_done) begin
          Stream2Mmap_13__state <= 2'b10;
        end 
      end 
      if(Stream2Mmap_13__state == 2'b10) begin
        if(Stream2Mmap_13__ap_done_global__q0) begin
          Stream2Mmap_13__state <= 2'b00;
        end 
      end 
    end
  end

  assign Stream2Mmap_13__ap_start = (Stream2Mmap_13__state == 2'b01);
  assign Stream2Mmap_14___n__q0 = n;
  assign Stream2Mmap_14___rmem14__q0 = rmem14;
  assign Stream2Mmap_14__ap_start_global__q0 = ap_start__q0;
  assign Stream2Mmap_14__is_done__q0 = (Stream2Mmap_14__state == 2'b10);
  assign Stream2Mmap_14__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Stream2Mmap_14__state <= 2'b00;
    end else begin
      if(Stream2Mmap_14__state == 2'b00) begin
        if(Stream2Mmap_14__ap_start_global__q0) begin
          Stream2Mmap_14__state <= 2'b01;
        end 
      end 
      if(Stream2Mmap_14__state == 2'b01) begin
        if(Stream2Mmap_14__ap_ready) begin
          if(Stream2Mmap_14__ap_done) begin
            Stream2Mmap_14__state <= 2'b10;
          end else begin
            Stream2Mmap_14__state <= 2'b11;
          end
        end 
      end 
      if(Stream2Mmap_14__state == 2'b11) begin
        if(Stream2Mmap_14__ap_done) begin
          Stream2Mmap_14__state <= 2'b10;
        end 
      end 
      if(Stream2Mmap_14__state == 2'b10) begin
        if(Stream2Mmap_14__ap_done_global__q0) begin
          Stream2Mmap_14__state <= 2'b00;
        end 
      end 
    end
  end

  assign Stream2Mmap_14__ap_start = (Stream2Mmap_14__state == 2'b01);
  assign Stream2Mmap_15___n__q0 = n;
  assign Stream2Mmap_15___rmem15__q0 = rmem15;
  assign Stream2Mmap_15__ap_start_global__q0 = ap_start__q0;
  assign Stream2Mmap_15__is_done__q0 = (Stream2Mmap_15__state == 2'b10);
  assign Stream2Mmap_15__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Stream2Mmap_15__state <= 2'b00;
    end else begin
      if(Stream2Mmap_15__state == 2'b00) begin
        if(Stream2Mmap_15__ap_start_global__q0) begin
          Stream2Mmap_15__state <= 2'b01;
        end 
      end 
      if(Stream2Mmap_15__state == 2'b01) begin
        if(Stream2Mmap_15__ap_ready) begin
          if(Stream2Mmap_15__ap_done) begin
            Stream2Mmap_15__state <= 2'b10;
          end else begin
            Stream2Mmap_15__state <= 2'b11;
          end
        end 
      end 
      if(Stream2Mmap_15__state == 2'b11) begin
        if(Stream2Mmap_15__ap_done) begin
          Stream2Mmap_15__state <= 2'b10;
        end 
      end 
      if(Stream2Mmap_15__state == 2'b10) begin
        if(Stream2Mmap_15__ap_done_global__q0) begin
          Stream2Mmap_15__state <= 2'b00;
        end 
      end 
    end
  end

  assign Stream2Mmap_15__ap_start = (Stream2Mmap_15__state == 2'b01);
  assign Stream2Mmap_16___n__q0 = n;
  assign Stream2Mmap_16___rmem16__q0 = rmem16;
  assign Stream2Mmap_16__ap_start_global__q0 = ap_start__q0;
  assign Stream2Mmap_16__is_done__q0 = (Stream2Mmap_16__state == 2'b10);
  assign Stream2Mmap_16__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Stream2Mmap_16__state <= 2'b00;
    end else begin
      if(Stream2Mmap_16__state == 2'b00) begin
        if(Stream2Mmap_16__ap_start_global__q0) begin
          Stream2Mmap_16__state <= 2'b01;
        end 
      end 
      if(Stream2Mmap_16__state == 2'b01) begin
        if(Stream2Mmap_16__ap_ready) begin
          if(Stream2Mmap_16__ap_done) begin
            Stream2Mmap_16__state <= 2'b10;
          end else begin
            Stream2Mmap_16__state <= 2'b11;
          end
        end 
      end 
      if(Stream2Mmap_16__state == 2'b11) begin
        if(Stream2Mmap_16__ap_done) begin
          Stream2Mmap_16__state <= 2'b10;
        end 
      end 
      if(Stream2Mmap_16__state == 2'b10) begin
        if(Stream2Mmap_16__ap_done_global__q0) begin
          Stream2Mmap_16__state <= 2'b00;
        end 
      end 
    end
  end

  assign Stream2Mmap_16__ap_start = (Stream2Mmap_16__state == 2'b01);
  assign Stream2Mmap_17___n__q0 = n;
  assign Stream2Mmap_17___rmem17__q0 = rmem17;
  assign Stream2Mmap_17__ap_start_global__q0 = ap_start__q0;
  assign Stream2Mmap_17__is_done__q0 = (Stream2Mmap_17__state == 2'b10);
  assign Stream2Mmap_17__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Stream2Mmap_17__state <= 2'b00;
    end else begin
      if(Stream2Mmap_17__state == 2'b00) begin
        if(Stream2Mmap_17__ap_start_global__q0) begin
          Stream2Mmap_17__state <= 2'b01;
        end 
      end 
      if(Stream2Mmap_17__state == 2'b01) begin
        if(Stream2Mmap_17__ap_ready) begin
          if(Stream2Mmap_17__ap_done) begin
            Stream2Mmap_17__state <= 2'b10;
          end else begin
            Stream2Mmap_17__state <= 2'b11;
          end
        end 
      end 
      if(Stream2Mmap_17__state == 2'b11) begin
        if(Stream2Mmap_17__ap_done) begin
          Stream2Mmap_17__state <= 2'b10;
        end 
      end 
      if(Stream2Mmap_17__state == 2'b10) begin
        if(Stream2Mmap_17__ap_done_global__q0) begin
          Stream2Mmap_17__state <= 2'b00;
        end 
      end 
    end
  end

  assign Stream2Mmap_17__ap_start = (Stream2Mmap_17__state == 2'b01);
  assign Stream2Mmap_18___n__q0 = n;
  assign Stream2Mmap_18___rmem18__q0 = rmem18;
  assign Stream2Mmap_18__ap_start_global__q0 = ap_start__q0;
  assign Stream2Mmap_18__is_done__q0 = (Stream2Mmap_18__state == 2'b10);
  assign Stream2Mmap_18__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Stream2Mmap_18__state <= 2'b00;
    end else begin
      if(Stream2Mmap_18__state == 2'b00) begin
        if(Stream2Mmap_18__ap_start_global__q0) begin
          Stream2Mmap_18__state <= 2'b01;
        end 
      end 
      if(Stream2Mmap_18__state == 2'b01) begin
        if(Stream2Mmap_18__ap_ready) begin
          if(Stream2Mmap_18__ap_done) begin
            Stream2Mmap_18__state <= 2'b10;
          end else begin
            Stream2Mmap_18__state <= 2'b11;
          end
        end 
      end 
      if(Stream2Mmap_18__state == 2'b11) begin
        if(Stream2Mmap_18__ap_done) begin
          Stream2Mmap_18__state <= 2'b10;
        end 
      end 
      if(Stream2Mmap_18__state == 2'b10) begin
        if(Stream2Mmap_18__ap_done_global__q0) begin
          Stream2Mmap_18__state <= 2'b00;
        end 
      end 
    end
  end

  assign Stream2Mmap_18__ap_start = (Stream2Mmap_18__state == 2'b01);
  assign Stream2Mmap_19___n__q0 = n;
  assign Stream2Mmap_19___rmem19__q0 = rmem19;
  assign Stream2Mmap_19__ap_start_global__q0 = ap_start__q0;
  assign Stream2Mmap_19__is_done__q0 = (Stream2Mmap_19__state == 2'b10);
  assign Stream2Mmap_19__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Stream2Mmap_19__state <= 2'b00;
    end else begin
      if(Stream2Mmap_19__state == 2'b00) begin
        if(Stream2Mmap_19__ap_start_global__q0) begin
          Stream2Mmap_19__state <= 2'b01;
        end 
      end 
      if(Stream2Mmap_19__state == 2'b01) begin
        if(Stream2Mmap_19__ap_ready) begin
          if(Stream2Mmap_19__ap_done) begin
            Stream2Mmap_19__state <= 2'b10;
          end else begin
            Stream2Mmap_19__state <= 2'b11;
          end
        end 
      end 
      if(Stream2Mmap_19__state == 2'b11) begin
        if(Stream2Mmap_19__ap_done) begin
          Stream2Mmap_19__state <= 2'b10;
        end 
      end 
      if(Stream2Mmap_19__state == 2'b10) begin
        if(Stream2Mmap_19__ap_done_global__q0) begin
          Stream2Mmap_19__state <= 2'b00;
        end 
      end 
    end
  end

  assign Stream2Mmap_19__ap_start = (Stream2Mmap_19__state == 2'b01);
  assign Stream2Mmap_20___n__q0 = n;
  assign Stream2Mmap_20___rmem20__q0 = rmem20;
  assign Stream2Mmap_20__ap_start_global__q0 = ap_start__q0;
  assign Stream2Mmap_20__is_done__q0 = (Stream2Mmap_20__state == 2'b10);
  assign Stream2Mmap_20__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Stream2Mmap_20__state <= 2'b00;
    end else begin
      if(Stream2Mmap_20__state == 2'b00) begin
        if(Stream2Mmap_20__ap_start_global__q0) begin
          Stream2Mmap_20__state <= 2'b01;
        end 
      end 
      if(Stream2Mmap_20__state == 2'b01) begin
        if(Stream2Mmap_20__ap_ready) begin
          if(Stream2Mmap_20__ap_done) begin
            Stream2Mmap_20__state <= 2'b10;
          end else begin
            Stream2Mmap_20__state <= 2'b11;
          end
        end 
      end 
      if(Stream2Mmap_20__state == 2'b11) begin
        if(Stream2Mmap_20__ap_done) begin
          Stream2Mmap_20__state <= 2'b10;
        end 
      end 
      if(Stream2Mmap_20__state == 2'b10) begin
        if(Stream2Mmap_20__ap_done_global__q0) begin
          Stream2Mmap_20__state <= 2'b00;
        end 
      end 
    end
  end

  assign Stream2Mmap_20__ap_start = (Stream2Mmap_20__state == 2'b01);
  assign Stream2Mmap_21___n__q0 = n;
  assign Stream2Mmap_21___rmem21__q0 = rmem21;
  assign Stream2Mmap_21__ap_start_global__q0 = ap_start__q0;
  assign Stream2Mmap_21__is_done__q0 = (Stream2Mmap_21__state == 2'b10);
  assign Stream2Mmap_21__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Stream2Mmap_21__state <= 2'b00;
    end else begin
      if(Stream2Mmap_21__state == 2'b00) begin
        if(Stream2Mmap_21__ap_start_global__q0) begin
          Stream2Mmap_21__state <= 2'b01;
        end 
      end 
      if(Stream2Mmap_21__state == 2'b01) begin
        if(Stream2Mmap_21__ap_ready) begin
          if(Stream2Mmap_21__ap_done) begin
            Stream2Mmap_21__state <= 2'b10;
          end else begin
            Stream2Mmap_21__state <= 2'b11;
          end
        end 
      end 
      if(Stream2Mmap_21__state == 2'b11) begin
        if(Stream2Mmap_21__ap_done) begin
          Stream2Mmap_21__state <= 2'b10;
        end 
      end 
      if(Stream2Mmap_21__state == 2'b10) begin
        if(Stream2Mmap_21__ap_done_global__q0) begin
          Stream2Mmap_21__state <= 2'b00;
        end 
      end 
    end
  end

  assign Stream2Mmap_21__ap_start = (Stream2Mmap_21__state == 2'b01);
  assign Stream2Mmap_22___n__q0 = n;
  assign Stream2Mmap_22___rmem22__q0 = rmem22;
  assign Stream2Mmap_22__ap_start_global__q0 = ap_start__q0;
  assign Stream2Mmap_22__is_done__q0 = (Stream2Mmap_22__state == 2'b10);
  assign Stream2Mmap_22__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Stream2Mmap_22__state <= 2'b00;
    end else begin
      if(Stream2Mmap_22__state == 2'b00) begin
        if(Stream2Mmap_22__ap_start_global__q0) begin
          Stream2Mmap_22__state <= 2'b01;
        end 
      end 
      if(Stream2Mmap_22__state == 2'b01) begin
        if(Stream2Mmap_22__ap_ready) begin
          if(Stream2Mmap_22__ap_done) begin
            Stream2Mmap_22__state <= 2'b10;
          end else begin
            Stream2Mmap_22__state <= 2'b11;
          end
        end 
      end 
      if(Stream2Mmap_22__state == 2'b11) begin
        if(Stream2Mmap_22__ap_done) begin
          Stream2Mmap_22__state <= 2'b10;
        end 
      end 
      if(Stream2Mmap_22__state == 2'b10) begin
        if(Stream2Mmap_22__ap_done_global__q0) begin
          Stream2Mmap_22__state <= 2'b00;
        end 
      end 
    end
  end

  assign Stream2Mmap_22__ap_start = (Stream2Mmap_22__state == 2'b01);
  assign Stream2Mmap_23___n__q0 = n;
  assign Stream2Mmap_23___rmem23__q0 = rmem23;
  assign Stream2Mmap_23__ap_start_global__q0 = ap_start__q0;
  assign Stream2Mmap_23__is_done__q0 = (Stream2Mmap_23__state == 2'b10);
  assign Stream2Mmap_23__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Stream2Mmap_23__state <= 2'b00;
    end else begin
      if(Stream2Mmap_23__state == 2'b00) begin
        if(Stream2Mmap_23__ap_start_global__q0) begin
          Stream2Mmap_23__state <= 2'b01;
        end 
      end 
      if(Stream2Mmap_23__state == 2'b01) begin
        if(Stream2Mmap_23__ap_ready) begin
          if(Stream2Mmap_23__ap_done) begin
            Stream2Mmap_23__state <= 2'b10;
          end else begin
            Stream2Mmap_23__state <= 2'b11;
          end
        end 
      end 
      if(Stream2Mmap_23__state == 2'b11) begin
        if(Stream2Mmap_23__ap_done) begin
          Stream2Mmap_23__state <= 2'b10;
        end 
      end 
      if(Stream2Mmap_23__state == 2'b10) begin
        if(Stream2Mmap_23__ap_done_global__q0) begin
          Stream2Mmap_23__state <= 2'b00;
        end 
      end 
    end
  end

  assign Stream2Mmap_23__ap_start = (Stream2Mmap_23__state == 2'b01);
  assign Stream2Mmap_24___n__q0 = n;
  assign Stream2Mmap_24___rmem24__q0 = rmem24;
  assign Stream2Mmap_24__ap_start_global__q0 = ap_start__q0;
  assign Stream2Mmap_24__is_done__q0 = (Stream2Mmap_24__state == 2'b10);
  assign Stream2Mmap_24__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Stream2Mmap_24__state <= 2'b00;
    end else begin
      if(Stream2Mmap_24__state == 2'b00) begin
        if(Stream2Mmap_24__ap_start_global__q0) begin
          Stream2Mmap_24__state <= 2'b01;
        end 
      end 
      if(Stream2Mmap_24__state == 2'b01) begin
        if(Stream2Mmap_24__ap_ready) begin
          if(Stream2Mmap_24__ap_done) begin
            Stream2Mmap_24__state <= 2'b10;
          end else begin
            Stream2Mmap_24__state <= 2'b11;
          end
        end 
      end 
      if(Stream2Mmap_24__state == 2'b11) begin
        if(Stream2Mmap_24__ap_done) begin
          Stream2Mmap_24__state <= 2'b10;
        end 
      end 
      if(Stream2Mmap_24__state == 2'b10) begin
        if(Stream2Mmap_24__ap_done_global__q0) begin
          Stream2Mmap_24__state <= 2'b00;
        end 
      end 
    end
  end

  assign Stream2Mmap_24__ap_start = (Stream2Mmap_24__state == 2'b01);
  assign Stream2Mmap_25___n__q0 = n;
  assign Stream2Mmap_25___rmem25__q0 = rmem25;
  assign Stream2Mmap_25__ap_start_global__q0 = ap_start__q0;
  assign Stream2Mmap_25__is_done__q0 = (Stream2Mmap_25__state == 2'b10);
  assign Stream2Mmap_25__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Stream2Mmap_25__state <= 2'b00;
    end else begin
      if(Stream2Mmap_25__state == 2'b00) begin
        if(Stream2Mmap_25__ap_start_global__q0) begin
          Stream2Mmap_25__state <= 2'b01;
        end 
      end 
      if(Stream2Mmap_25__state == 2'b01) begin
        if(Stream2Mmap_25__ap_ready) begin
          if(Stream2Mmap_25__ap_done) begin
            Stream2Mmap_25__state <= 2'b10;
          end else begin
            Stream2Mmap_25__state <= 2'b11;
          end
        end 
      end 
      if(Stream2Mmap_25__state == 2'b11) begin
        if(Stream2Mmap_25__ap_done) begin
          Stream2Mmap_25__state <= 2'b10;
        end 
      end 
      if(Stream2Mmap_25__state == 2'b10) begin
        if(Stream2Mmap_25__ap_done_global__q0) begin
          Stream2Mmap_25__state <= 2'b00;
        end 
      end 
    end
  end

  assign Stream2Mmap_25__ap_start = (Stream2Mmap_25__state == 2'b01);
  assign Stream2Mmap_26___n__q0 = n;
  assign Stream2Mmap_26___rmem26__q0 = rmem26;
  assign Stream2Mmap_26__ap_start_global__q0 = ap_start__q0;
  assign Stream2Mmap_26__is_done__q0 = (Stream2Mmap_26__state == 2'b10);
  assign Stream2Mmap_26__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Stream2Mmap_26__state <= 2'b00;
    end else begin
      if(Stream2Mmap_26__state == 2'b00) begin
        if(Stream2Mmap_26__ap_start_global__q0) begin
          Stream2Mmap_26__state <= 2'b01;
        end 
      end 
      if(Stream2Mmap_26__state == 2'b01) begin
        if(Stream2Mmap_26__ap_ready) begin
          if(Stream2Mmap_26__ap_done) begin
            Stream2Mmap_26__state <= 2'b10;
          end else begin
            Stream2Mmap_26__state <= 2'b11;
          end
        end 
      end 
      if(Stream2Mmap_26__state == 2'b11) begin
        if(Stream2Mmap_26__ap_done) begin
          Stream2Mmap_26__state <= 2'b10;
        end 
      end 
      if(Stream2Mmap_26__state == 2'b10) begin
        if(Stream2Mmap_26__ap_done_global__q0) begin
          Stream2Mmap_26__state <= 2'b00;
        end 
      end 
    end
  end

  assign Stream2Mmap_26__ap_start = (Stream2Mmap_26__state == 2'b01);
  assign yshift_0___n__q0 = n;
  assign yshift_0__ap_start_global__q0 = ap_start__q0;
  assign yshift_0__is_done__q0 = (yshift_0__state == 2'b10);
  assign yshift_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yshift_0__state <= 2'b00;
    end else begin
      if(yshift_0__state == 2'b00) begin
        if(yshift_0__ap_start_global__q0) begin
          yshift_0__state <= 2'b01;
        end 
      end 
      if(yshift_0__state == 2'b01) begin
        if(yshift_0__ap_ready) begin
          if(yshift_0__ap_done) begin
            yshift_0__state <= 2'b10;
          end else begin
            yshift_0__state <= 2'b11;
          end
        end 
      end 
      if(yshift_0__state == 2'b11) begin
        if(yshift_0__ap_done) begin
          yshift_0__state <= 2'b10;
        end 
      end 
      if(yshift_0__state == 2'b10) begin
        if(yshift_0__ap_done_global__q0) begin
          yshift_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign yshift_0__ap_start = (yshift_0__state == 2'b01);
  assign yshift_1___n__q0 = n;
  assign yshift_1__ap_start_global__q0 = ap_start__q0;
  assign yshift_1__is_done__q0 = (yshift_1__state == 2'b10);
  assign yshift_1__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yshift_1__state <= 2'b00;
    end else begin
      if(yshift_1__state == 2'b00) begin
        if(yshift_1__ap_start_global__q0) begin
          yshift_1__state <= 2'b01;
        end 
      end 
      if(yshift_1__state == 2'b01) begin
        if(yshift_1__ap_ready) begin
          if(yshift_1__ap_done) begin
            yshift_1__state <= 2'b10;
          end else begin
            yshift_1__state <= 2'b11;
          end
        end 
      end 
      if(yshift_1__state == 2'b11) begin
        if(yshift_1__ap_done) begin
          yshift_1__state <= 2'b10;
        end 
      end 
      if(yshift_1__state == 2'b10) begin
        if(yshift_1__ap_done_global__q0) begin
          yshift_1__state <= 2'b00;
        end 
      end 
    end
  end

  assign yshift_1__ap_start = (yshift_1__state == 2'b01);
  assign yshift_2___n__q0 = n;
  assign yshift_2__ap_start_global__q0 = ap_start__q0;
  assign yshift_2__is_done__q0 = (yshift_2__state == 2'b10);
  assign yshift_2__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yshift_2__state <= 2'b00;
    end else begin
      if(yshift_2__state == 2'b00) begin
        if(yshift_2__ap_start_global__q0) begin
          yshift_2__state <= 2'b01;
        end 
      end 
      if(yshift_2__state == 2'b01) begin
        if(yshift_2__ap_ready) begin
          if(yshift_2__ap_done) begin
            yshift_2__state <= 2'b10;
          end else begin
            yshift_2__state <= 2'b11;
          end
        end 
      end 
      if(yshift_2__state == 2'b11) begin
        if(yshift_2__ap_done) begin
          yshift_2__state <= 2'b10;
        end 
      end 
      if(yshift_2__state == 2'b10) begin
        if(yshift_2__ap_done_global__q0) begin
          yshift_2__state <= 2'b00;
        end 
      end 
    end
  end

  assign yshift_2__ap_start = (yshift_2__state == 2'b01);
  assign yshift_3___n__q0 = n;
  assign yshift_3__ap_start_global__q0 = ap_start__q0;
  assign yshift_3__is_done__q0 = (yshift_3__state == 2'b10);
  assign yshift_3__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yshift_3__state <= 2'b00;
    end else begin
      if(yshift_3__state == 2'b00) begin
        if(yshift_3__ap_start_global__q0) begin
          yshift_3__state <= 2'b01;
        end 
      end 
      if(yshift_3__state == 2'b01) begin
        if(yshift_3__ap_ready) begin
          if(yshift_3__ap_done) begin
            yshift_3__state <= 2'b10;
          end else begin
            yshift_3__state <= 2'b11;
          end
        end 
      end 
      if(yshift_3__state == 2'b11) begin
        if(yshift_3__ap_done) begin
          yshift_3__state <= 2'b10;
        end 
      end 
      if(yshift_3__state == 2'b10) begin
        if(yshift_3__ap_done_global__q0) begin
          yshift_3__state <= 2'b00;
        end 
      end 
    end
  end

  assign yshift_3__ap_start = (yshift_3__state == 2'b01);
  assign yshift_4___n__q0 = n;
  assign yshift_4__ap_start_global__q0 = ap_start__q0;
  assign yshift_4__is_done__q0 = (yshift_4__state == 2'b10);
  assign yshift_4__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yshift_4__state <= 2'b00;
    end else begin
      if(yshift_4__state == 2'b00) begin
        if(yshift_4__ap_start_global__q0) begin
          yshift_4__state <= 2'b01;
        end 
      end 
      if(yshift_4__state == 2'b01) begin
        if(yshift_4__ap_ready) begin
          if(yshift_4__ap_done) begin
            yshift_4__state <= 2'b10;
          end else begin
            yshift_4__state <= 2'b11;
          end
        end 
      end 
      if(yshift_4__state == 2'b11) begin
        if(yshift_4__ap_done) begin
          yshift_4__state <= 2'b10;
        end 
      end 
      if(yshift_4__state == 2'b10) begin
        if(yshift_4__ap_done_global__q0) begin
          yshift_4__state <= 2'b00;
        end 
      end 
    end
  end

  assign yshift_4__ap_start = (yshift_4__state == 2'b01);
  assign yshift_5___n__q0 = n;
  assign yshift_5__ap_start_global__q0 = ap_start__q0;
  assign yshift_5__is_done__q0 = (yshift_5__state == 2'b10);
  assign yshift_5__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yshift_5__state <= 2'b00;
    end else begin
      if(yshift_5__state == 2'b00) begin
        if(yshift_5__ap_start_global__q0) begin
          yshift_5__state <= 2'b01;
        end 
      end 
      if(yshift_5__state == 2'b01) begin
        if(yshift_5__ap_ready) begin
          if(yshift_5__ap_done) begin
            yshift_5__state <= 2'b10;
          end else begin
            yshift_5__state <= 2'b11;
          end
        end 
      end 
      if(yshift_5__state == 2'b11) begin
        if(yshift_5__ap_done) begin
          yshift_5__state <= 2'b10;
        end 
      end 
      if(yshift_5__state == 2'b10) begin
        if(yshift_5__ap_done_global__q0) begin
          yshift_5__state <= 2'b00;
        end 
      end 
    end
  end

  assign yshift_5__ap_start = (yshift_5__state == 2'b01);
  assign yshift_6___n__q0 = n;
  assign yshift_6__ap_start_global__q0 = ap_start__q0;
  assign yshift_6__is_done__q0 = (yshift_6__state == 2'b10);
  assign yshift_6__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yshift_6__state <= 2'b00;
    end else begin
      if(yshift_6__state == 2'b00) begin
        if(yshift_6__ap_start_global__q0) begin
          yshift_6__state <= 2'b01;
        end 
      end 
      if(yshift_6__state == 2'b01) begin
        if(yshift_6__ap_ready) begin
          if(yshift_6__ap_done) begin
            yshift_6__state <= 2'b10;
          end else begin
            yshift_6__state <= 2'b11;
          end
        end 
      end 
      if(yshift_6__state == 2'b11) begin
        if(yshift_6__ap_done) begin
          yshift_6__state <= 2'b10;
        end 
      end 
      if(yshift_6__state == 2'b10) begin
        if(yshift_6__ap_done_global__q0) begin
          yshift_6__state <= 2'b00;
        end 
      end 
    end
  end

  assign yshift_6__ap_start = (yshift_6__state == 2'b01);
  assign yshift_7___n__q0 = n;
  assign yshift_7__ap_start_global__q0 = ap_start__q0;
  assign yshift_7__is_done__q0 = (yshift_7__state == 2'b10);
  assign yshift_7__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yshift_7__state <= 2'b00;
    end else begin
      if(yshift_7__state == 2'b00) begin
        if(yshift_7__ap_start_global__q0) begin
          yshift_7__state <= 2'b01;
        end 
      end 
      if(yshift_7__state == 2'b01) begin
        if(yshift_7__ap_ready) begin
          if(yshift_7__ap_done) begin
            yshift_7__state <= 2'b10;
          end else begin
            yshift_7__state <= 2'b11;
          end
        end 
      end 
      if(yshift_7__state == 2'b11) begin
        if(yshift_7__ap_done) begin
          yshift_7__state <= 2'b10;
        end 
      end 
      if(yshift_7__state == 2'b10) begin
        if(yshift_7__ap_done_global__q0) begin
          yshift_7__state <= 2'b00;
        end 
      end 
    end
  end

  assign yshift_7__ap_start = (yshift_7__state == 2'b01);
  assign yshift_8___n__q0 = n;
  assign yshift_8__ap_start_global__q0 = ap_start__q0;
  assign yshift_8__is_done__q0 = (yshift_8__state == 2'b10);
  assign yshift_8__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yshift_8__state <= 2'b00;
    end else begin
      if(yshift_8__state == 2'b00) begin
        if(yshift_8__ap_start_global__q0) begin
          yshift_8__state <= 2'b01;
        end 
      end 
      if(yshift_8__state == 2'b01) begin
        if(yshift_8__ap_ready) begin
          if(yshift_8__ap_done) begin
            yshift_8__state <= 2'b10;
          end else begin
            yshift_8__state <= 2'b11;
          end
        end 
      end 
      if(yshift_8__state == 2'b11) begin
        if(yshift_8__ap_done) begin
          yshift_8__state <= 2'b10;
        end 
      end 
      if(yshift_8__state == 2'b10) begin
        if(yshift_8__ap_done_global__q0) begin
          yshift_8__state <= 2'b00;
        end 
      end 
    end
  end

  assign yshift_8__ap_start = (yshift_8__state == 2'b01);
  assign yshift_9___n__q0 = n;
  assign yshift_9__ap_start_global__q0 = ap_start__q0;
  assign yshift_9__is_done__q0 = (yshift_9__state == 2'b10);
  assign yshift_9__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yshift_9__state <= 2'b00;
    end else begin
      if(yshift_9__state == 2'b00) begin
        if(yshift_9__ap_start_global__q0) begin
          yshift_9__state <= 2'b01;
        end 
      end 
      if(yshift_9__state == 2'b01) begin
        if(yshift_9__ap_ready) begin
          if(yshift_9__ap_done) begin
            yshift_9__state <= 2'b10;
          end else begin
            yshift_9__state <= 2'b11;
          end
        end 
      end 
      if(yshift_9__state == 2'b11) begin
        if(yshift_9__ap_done) begin
          yshift_9__state <= 2'b10;
        end 
      end 
      if(yshift_9__state == 2'b10) begin
        if(yshift_9__ap_done_global__q0) begin
          yshift_9__state <= 2'b00;
        end 
      end 
    end
  end

  assign yshift_9__ap_start = (yshift_9__state == 2'b01);
  assign yshift_10___n__q0 = n;
  assign yshift_10__ap_start_global__q0 = ap_start__q0;
  assign yshift_10__is_done__q0 = (yshift_10__state == 2'b10);
  assign yshift_10__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yshift_10__state <= 2'b00;
    end else begin
      if(yshift_10__state == 2'b00) begin
        if(yshift_10__ap_start_global__q0) begin
          yshift_10__state <= 2'b01;
        end 
      end 
      if(yshift_10__state == 2'b01) begin
        if(yshift_10__ap_ready) begin
          if(yshift_10__ap_done) begin
            yshift_10__state <= 2'b10;
          end else begin
            yshift_10__state <= 2'b11;
          end
        end 
      end 
      if(yshift_10__state == 2'b11) begin
        if(yshift_10__ap_done) begin
          yshift_10__state <= 2'b10;
        end 
      end 
      if(yshift_10__state == 2'b10) begin
        if(yshift_10__ap_done_global__q0) begin
          yshift_10__state <= 2'b00;
        end 
      end 
    end
  end

  assign yshift_10__ap_start = (yshift_10__state == 2'b01);
  assign yshift_11___n__q0 = n;
  assign yshift_11__ap_start_global__q0 = ap_start__q0;
  assign yshift_11__is_done__q0 = (yshift_11__state == 2'b10);
  assign yshift_11__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yshift_11__state <= 2'b00;
    end else begin
      if(yshift_11__state == 2'b00) begin
        if(yshift_11__ap_start_global__q0) begin
          yshift_11__state <= 2'b01;
        end 
      end 
      if(yshift_11__state == 2'b01) begin
        if(yshift_11__ap_ready) begin
          if(yshift_11__ap_done) begin
            yshift_11__state <= 2'b10;
          end else begin
            yshift_11__state <= 2'b11;
          end
        end 
      end 
      if(yshift_11__state == 2'b11) begin
        if(yshift_11__ap_done) begin
          yshift_11__state <= 2'b10;
        end 
      end 
      if(yshift_11__state == 2'b10) begin
        if(yshift_11__ap_done_global__q0) begin
          yshift_11__state <= 2'b00;
        end 
      end 
    end
  end

  assign yshift_11__ap_start = (yshift_11__state == 2'b01);
  assign yshift_12___n__q0 = n;
  assign yshift_12__ap_start_global__q0 = ap_start__q0;
  assign yshift_12__is_done__q0 = (yshift_12__state == 2'b10);
  assign yshift_12__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yshift_12__state <= 2'b00;
    end else begin
      if(yshift_12__state == 2'b00) begin
        if(yshift_12__ap_start_global__q0) begin
          yshift_12__state <= 2'b01;
        end 
      end 
      if(yshift_12__state == 2'b01) begin
        if(yshift_12__ap_ready) begin
          if(yshift_12__ap_done) begin
            yshift_12__state <= 2'b10;
          end else begin
            yshift_12__state <= 2'b11;
          end
        end 
      end 
      if(yshift_12__state == 2'b11) begin
        if(yshift_12__ap_done) begin
          yshift_12__state <= 2'b10;
        end 
      end 
      if(yshift_12__state == 2'b10) begin
        if(yshift_12__ap_done_global__q0) begin
          yshift_12__state <= 2'b00;
        end 
      end 
    end
  end

  assign yshift_12__ap_start = (yshift_12__state == 2'b01);
  assign yshift_13___n__q0 = n;
  assign yshift_13__ap_start_global__q0 = ap_start__q0;
  assign yshift_13__is_done__q0 = (yshift_13__state == 2'b10);
  assign yshift_13__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yshift_13__state <= 2'b00;
    end else begin
      if(yshift_13__state == 2'b00) begin
        if(yshift_13__ap_start_global__q0) begin
          yshift_13__state <= 2'b01;
        end 
      end 
      if(yshift_13__state == 2'b01) begin
        if(yshift_13__ap_ready) begin
          if(yshift_13__ap_done) begin
            yshift_13__state <= 2'b10;
          end else begin
            yshift_13__state <= 2'b11;
          end
        end 
      end 
      if(yshift_13__state == 2'b11) begin
        if(yshift_13__ap_done) begin
          yshift_13__state <= 2'b10;
        end 
      end 
      if(yshift_13__state == 2'b10) begin
        if(yshift_13__ap_done_global__q0) begin
          yshift_13__state <= 2'b00;
        end 
      end 
    end
  end

  assign yshift_13__ap_start = (yshift_13__state == 2'b01);
  assign yshift_14___n__q0 = n;
  assign yshift_14__ap_start_global__q0 = ap_start__q0;
  assign yshift_14__is_done__q0 = (yshift_14__state == 2'b10);
  assign yshift_14__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yshift_14__state <= 2'b00;
    end else begin
      if(yshift_14__state == 2'b00) begin
        if(yshift_14__ap_start_global__q0) begin
          yshift_14__state <= 2'b01;
        end 
      end 
      if(yshift_14__state == 2'b01) begin
        if(yshift_14__ap_ready) begin
          if(yshift_14__ap_done) begin
            yshift_14__state <= 2'b10;
          end else begin
            yshift_14__state <= 2'b11;
          end
        end 
      end 
      if(yshift_14__state == 2'b11) begin
        if(yshift_14__ap_done) begin
          yshift_14__state <= 2'b10;
        end 
      end 
      if(yshift_14__state == 2'b10) begin
        if(yshift_14__ap_done_global__q0) begin
          yshift_14__state <= 2'b00;
        end 
      end 
    end
  end

  assign yshift_14__ap_start = (yshift_14__state == 2'b01);
  assign yshift_15___n__q0 = n;
  assign yshift_15__ap_start_global__q0 = ap_start__q0;
  assign yshift_15__is_done__q0 = (yshift_15__state == 2'b10);
  assign yshift_15__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yshift_15__state <= 2'b00;
    end else begin
      if(yshift_15__state == 2'b00) begin
        if(yshift_15__ap_start_global__q0) begin
          yshift_15__state <= 2'b01;
        end 
      end 
      if(yshift_15__state == 2'b01) begin
        if(yshift_15__ap_ready) begin
          if(yshift_15__ap_done) begin
            yshift_15__state <= 2'b10;
          end else begin
            yshift_15__state <= 2'b11;
          end
        end 
      end 
      if(yshift_15__state == 2'b11) begin
        if(yshift_15__ap_done) begin
          yshift_15__state <= 2'b10;
        end 
      end 
      if(yshift_15__state == 2'b10) begin
        if(yshift_15__ap_done_global__q0) begin
          yshift_15__state <= 2'b00;
        end 
      end 
    end
  end

  assign yshift_15__ap_start = (yshift_15__state == 2'b01);
  assign yshift_16___n__q0 = n;
  assign yshift_16__ap_start_global__q0 = ap_start__q0;
  assign yshift_16__is_done__q0 = (yshift_16__state == 2'b10);
  assign yshift_16__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yshift_16__state <= 2'b00;
    end else begin
      if(yshift_16__state == 2'b00) begin
        if(yshift_16__ap_start_global__q0) begin
          yshift_16__state <= 2'b01;
        end 
      end 
      if(yshift_16__state == 2'b01) begin
        if(yshift_16__ap_ready) begin
          if(yshift_16__ap_done) begin
            yshift_16__state <= 2'b10;
          end else begin
            yshift_16__state <= 2'b11;
          end
        end 
      end 
      if(yshift_16__state == 2'b11) begin
        if(yshift_16__ap_done) begin
          yshift_16__state <= 2'b10;
        end 
      end 
      if(yshift_16__state == 2'b10) begin
        if(yshift_16__ap_done_global__q0) begin
          yshift_16__state <= 2'b00;
        end 
      end 
    end
  end

  assign yshift_16__ap_start = (yshift_16__state == 2'b01);
  assign yshift_17___n__q0 = n;
  assign yshift_17__ap_start_global__q0 = ap_start__q0;
  assign yshift_17__is_done__q0 = (yshift_17__state == 2'b10);
  assign yshift_17__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yshift_17__state <= 2'b00;
    end else begin
      if(yshift_17__state == 2'b00) begin
        if(yshift_17__ap_start_global__q0) begin
          yshift_17__state <= 2'b01;
        end 
      end 
      if(yshift_17__state == 2'b01) begin
        if(yshift_17__ap_ready) begin
          if(yshift_17__ap_done) begin
            yshift_17__state <= 2'b10;
          end else begin
            yshift_17__state <= 2'b11;
          end
        end 
      end 
      if(yshift_17__state == 2'b11) begin
        if(yshift_17__ap_done) begin
          yshift_17__state <= 2'b10;
        end 
      end 
      if(yshift_17__state == 2'b10) begin
        if(yshift_17__ap_done_global__q0) begin
          yshift_17__state <= 2'b00;
        end 
      end 
    end
  end

  assign yshift_17__ap_start = (yshift_17__state == 2'b01);
  assign yshift_18___n__q0 = n;
  assign yshift_18__ap_start_global__q0 = ap_start__q0;
  assign yshift_18__is_done__q0 = (yshift_18__state == 2'b10);
  assign yshift_18__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yshift_18__state <= 2'b00;
    end else begin
      if(yshift_18__state == 2'b00) begin
        if(yshift_18__ap_start_global__q0) begin
          yshift_18__state <= 2'b01;
        end 
      end 
      if(yshift_18__state == 2'b01) begin
        if(yshift_18__ap_ready) begin
          if(yshift_18__ap_done) begin
            yshift_18__state <= 2'b10;
          end else begin
            yshift_18__state <= 2'b11;
          end
        end 
      end 
      if(yshift_18__state == 2'b11) begin
        if(yshift_18__ap_done) begin
          yshift_18__state <= 2'b10;
        end 
      end 
      if(yshift_18__state == 2'b10) begin
        if(yshift_18__ap_done_global__q0) begin
          yshift_18__state <= 2'b00;
        end 
      end 
    end
  end

  assign yshift_18__ap_start = (yshift_18__state == 2'b01);
  assign yshift_19___n__q0 = n;
  assign yshift_19__ap_start_global__q0 = ap_start__q0;
  assign yshift_19__is_done__q0 = (yshift_19__state == 2'b10);
  assign yshift_19__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yshift_19__state <= 2'b00;
    end else begin
      if(yshift_19__state == 2'b00) begin
        if(yshift_19__ap_start_global__q0) begin
          yshift_19__state <= 2'b01;
        end 
      end 
      if(yshift_19__state == 2'b01) begin
        if(yshift_19__ap_ready) begin
          if(yshift_19__ap_done) begin
            yshift_19__state <= 2'b10;
          end else begin
            yshift_19__state <= 2'b11;
          end
        end 
      end 
      if(yshift_19__state == 2'b11) begin
        if(yshift_19__ap_done) begin
          yshift_19__state <= 2'b10;
        end 
      end 
      if(yshift_19__state == 2'b10) begin
        if(yshift_19__ap_done_global__q0) begin
          yshift_19__state <= 2'b00;
        end 
      end 
    end
  end

  assign yshift_19__ap_start = (yshift_19__state == 2'b01);
  assign yshift_20___n__q0 = n;
  assign yshift_20__ap_start_global__q0 = ap_start__q0;
  assign yshift_20__is_done__q0 = (yshift_20__state == 2'b10);
  assign yshift_20__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yshift_20__state <= 2'b00;
    end else begin
      if(yshift_20__state == 2'b00) begin
        if(yshift_20__ap_start_global__q0) begin
          yshift_20__state <= 2'b01;
        end 
      end 
      if(yshift_20__state == 2'b01) begin
        if(yshift_20__ap_ready) begin
          if(yshift_20__ap_done) begin
            yshift_20__state <= 2'b10;
          end else begin
            yshift_20__state <= 2'b11;
          end
        end 
      end 
      if(yshift_20__state == 2'b11) begin
        if(yshift_20__ap_done) begin
          yshift_20__state <= 2'b10;
        end 
      end 
      if(yshift_20__state == 2'b10) begin
        if(yshift_20__ap_done_global__q0) begin
          yshift_20__state <= 2'b00;
        end 
      end 
    end
  end

  assign yshift_20__ap_start = (yshift_20__state == 2'b01);
  assign yshift_21___n__q0 = n;
  assign yshift_21__ap_start_global__q0 = ap_start__q0;
  assign yshift_21__is_done__q0 = (yshift_21__state == 2'b10);
  assign yshift_21__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yshift_21__state <= 2'b00;
    end else begin
      if(yshift_21__state == 2'b00) begin
        if(yshift_21__ap_start_global__q0) begin
          yshift_21__state <= 2'b01;
        end 
      end 
      if(yshift_21__state == 2'b01) begin
        if(yshift_21__ap_ready) begin
          if(yshift_21__ap_done) begin
            yshift_21__state <= 2'b10;
          end else begin
            yshift_21__state <= 2'b11;
          end
        end 
      end 
      if(yshift_21__state == 2'b11) begin
        if(yshift_21__ap_done) begin
          yshift_21__state <= 2'b10;
        end 
      end 
      if(yshift_21__state == 2'b10) begin
        if(yshift_21__ap_done_global__q0) begin
          yshift_21__state <= 2'b00;
        end 
      end 
    end
  end

  assign yshift_21__ap_start = (yshift_21__state == 2'b01);
  assign yshift_22___n__q0 = n;
  assign yshift_22__ap_start_global__q0 = ap_start__q0;
  assign yshift_22__is_done__q0 = (yshift_22__state == 2'b10);
  assign yshift_22__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yshift_22__state <= 2'b00;
    end else begin
      if(yshift_22__state == 2'b00) begin
        if(yshift_22__ap_start_global__q0) begin
          yshift_22__state <= 2'b01;
        end 
      end 
      if(yshift_22__state == 2'b01) begin
        if(yshift_22__ap_ready) begin
          if(yshift_22__ap_done) begin
            yshift_22__state <= 2'b10;
          end else begin
            yshift_22__state <= 2'b11;
          end
        end 
      end 
      if(yshift_22__state == 2'b11) begin
        if(yshift_22__ap_done) begin
          yshift_22__state <= 2'b10;
        end 
      end 
      if(yshift_22__state == 2'b10) begin
        if(yshift_22__ap_done_global__q0) begin
          yshift_22__state <= 2'b00;
        end 
      end 
    end
  end

  assign yshift_22__ap_start = (yshift_22__state == 2'b01);
  assign yshift_23___n__q0 = n;
  assign yshift_23__ap_start_global__q0 = ap_start__q0;
  assign yshift_23__is_done__q0 = (yshift_23__state == 2'b10);
  assign yshift_23__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yshift_23__state <= 2'b00;
    end else begin
      if(yshift_23__state == 2'b00) begin
        if(yshift_23__ap_start_global__q0) begin
          yshift_23__state <= 2'b01;
        end 
      end 
      if(yshift_23__state == 2'b01) begin
        if(yshift_23__ap_ready) begin
          if(yshift_23__ap_done) begin
            yshift_23__state <= 2'b10;
          end else begin
            yshift_23__state <= 2'b11;
          end
        end 
      end 
      if(yshift_23__state == 2'b11) begin
        if(yshift_23__ap_done) begin
          yshift_23__state <= 2'b10;
        end 
      end 
      if(yshift_23__state == 2'b10) begin
        if(yshift_23__ap_done_global__q0) begin
          yshift_23__state <= 2'b00;
        end 
      end 
    end
  end

  assign yshift_23__ap_start = (yshift_23__state == 2'b01);
  assign yshift_24___n__q0 = n;
  assign yshift_24__ap_start_global__q0 = ap_start__q0;
  assign yshift_24__is_done__q0 = (yshift_24__state == 2'b10);
  assign yshift_24__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yshift_24__state <= 2'b00;
    end else begin
      if(yshift_24__state == 2'b00) begin
        if(yshift_24__ap_start_global__q0) begin
          yshift_24__state <= 2'b01;
        end 
      end 
      if(yshift_24__state == 2'b01) begin
        if(yshift_24__ap_ready) begin
          if(yshift_24__ap_done) begin
            yshift_24__state <= 2'b10;
          end else begin
            yshift_24__state <= 2'b11;
          end
        end 
      end 
      if(yshift_24__state == 2'b11) begin
        if(yshift_24__ap_done) begin
          yshift_24__state <= 2'b10;
        end 
      end 
      if(yshift_24__state == 2'b10) begin
        if(yshift_24__ap_done_global__q0) begin
          yshift_24__state <= 2'b00;
        end 
      end 
    end
  end

  assign yshift_24__ap_start = (yshift_24__state == 2'b01);
  assign yshift_25___n__q0 = n;
  assign yshift_25__ap_start_global__q0 = ap_start__q0;
  assign yshift_25__is_done__q0 = (yshift_25__state == 2'b10);
  assign yshift_25__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yshift_25__state <= 2'b00;
    end else begin
      if(yshift_25__state == 2'b00) begin
        if(yshift_25__ap_start_global__q0) begin
          yshift_25__state <= 2'b01;
        end 
      end 
      if(yshift_25__state == 2'b01) begin
        if(yshift_25__ap_ready) begin
          if(yshift_25__ap_done) begin
            yshift_25__state <= 2'b10;
          end else begin
            yshift_25__state <= 2'b11;
          end
        end 
      end 
      if(yshift_25__state == 2'b11) begin
        if(yshift_25__ap_done) begin
          yshift_25__state <= 2'b10;
        end 
      end 
      if(yshift_25__state == 2'b10) begin
        if(yshift_25__ap_done_global__q0) begin
          yshift_25__state <= 2'b00;
        end 
      end 
    end
  end

  assign yshift_25__ap_start = (yshift_25__state == 2'b01);
  assign yshift_26___n__q0 = n;
  assign yshift_26__ap_start_global__q0 = ap_start__q0;
  assign yshift_26__is_done__q0 = (yshift_26__state == 2'b10);
  assign yshift_26__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      yshift_26__state <= 2'b00;
    end else begin
      if(yshift_26__state == 2'b00) begin
        if(yshift_26__ap_start_global__q0) begin
          yshift_26__state <= 2'b01;
        end 
      end 
      if(yshift_26__state == 2'b01) begin
        if(yshift_26__ap_ready) begin
          if(yshift_26__ap_done) begin
            yshift_26__state <= 2'b10;
          end else begin
            yshift_26__state <= 2'b11;
          end
        end 
      end 
      if(yshift_26__state == 2'b11) begin
        if(yshift_26__ap_done) begin
          yshift_26__state <= 2'b10;
        end 
      end 
      if(yshift_26__state == 2'b10) begin
        if(yshift_26__ap_done_global__q0) begin
          yshift_26__state <= 2'b00;
        end 
      end 
    end
  end

  assign yshift_26__ap_start = (yshift_26__state == 2'b01);

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      tapa_state <= 2'b00;
    end else begin
      case(tapa_state)
        2'b00: begin
          if(ap_start__q0) begin
            tapa_state <= 2'b01;
          end 
        end
        2'b01: begin
          if(Mmap2Stream_0__is_done__q0 && Mmap2Stream_1__is_done__q0 && Mmap2Stream_2__is_done__q0 && Mmap2Stream_3__is_done__q0 && Mmap2Stream_4__is_done__q0 && Mmap2Stream_5__is_done__q0 && Mmap2Stream_6__is_done__q0 && Mmap2Stream_7__is_done__q0 && Mmap2Stream_8__is_done__q0 && Mmap2Stream_9__is_done__q0 && Mmap2Stream_10__is_done__q0 && Mmap2Stream_11__is_done__q0 && Mmap2Stream_12__is_done__q0 && Mmap2Stream_13__is_done__q0 && Mmap2Stream_14__is_done__q0 && Mmap2Stream_15__is_done__q0 && Mmap2Stream_16__is_done__q0 && Mmap2Stream_17__is_done__q0 && Mmap2Stream_18__is_done__q0 && Mmap2Stream_19__is_done__q0 && Mmap2Stream_20__is_done__q0 && Mmap2Stream_21__is_done__q0 && Mmap2Stream_22__is_done__q0 && Mmap2Stream_23__is_done__q0 && Mmap2Stream_24__is_done__q0 && Mmap2Stream_25__is_done__q0 && Mmap2Stream_26__is_done__q0 && Stream2Mmap_0__is_done__q0 && Stream2Mmap_1__is_done__q0 && Stream2Mmap_2__is_done__q0 && Stream2Mmap_3__is_done__q0 && Stream2Mmap_4__is_done__q0 && Stream2Mmap_5__is_done__q0 && Stream2Mmap_6__is_done__q0 && Stream2Mmap_7__is_done__q0 && Stream2Mmap_8__is_done__q0 && Stream2Mmap_9__is_done__q0 && Stream2Mmap_10__is_done__q0 && Stream2Mmap_11__is_done__q0 && Stream2Mmap_12__is_done__q0 && Stream2Mmap_13__is_done__q0 && Stream2Mmap_14__is_done__q0 && Stream2Mmap_15__is_done__q0 && Stream2Mmap_16__is_done__q0 && Stream2Mmap_17__is_done__q0 && Stream2Mmap_18__is_done__q0 && Stream2Mmap_19__is_done__q0 && Stream2Mmap_20__is_done__q0 && Stream2Mmap_21__is_done__q0 && Stream2Mmap_22__is_done__q0 && Stream2Mmap_23__is_done__q0 && Stream2Mmap_24__is_done__q0 && Stream2Mmap_25__is_done__q0 && Stream2Mmap_26__is_done__q0 && yshift_0__is_done__q0 && yshift_1__is_done__q0 && yshift_2__is_done__q0 && yshift_3__is_done__q0 && yshift_4__is_done__q0 && yshift_5__is_done__q0 && yshift_6__is_done__q0 && yshift_7__is_done__q0 && yshift_8__is_done__q0 && yshift_9__is_done__q0 && yshift_10__is_done__q0 && yshift_11__is_done__q0 && yshift_12__is_done__q0 && yshift_13__is_done__q0 && yshift_14__is_done__q0 && yshift_15__is_done__q0 && yshift_16__is_done__q0 && yshift_17__is_done__q0 && yshift_18__is_done__q0 && yshift_19__is_done__q0 && yshift_20__is_done__q0 && yshift_21__is_done__q0 && yshift_22__is_done__q0 && yshift_23__is_done__q0 && yshift_24__is_done__q0 && yshift_25__is_done__q0 && yshift_26__is_done__q0) begin
            tapa_state <= 2'b10;
          end 
        end
        2'b10: begin
          tapa_state <= 2'b00;
          countdown <= 1'd0;
        end
        2'b11: begin
          if(countdown == 1'd0) begin
            tapa_state <= 2'b00;
          end else begin
            countdown <= (countdown - 1'd1);
          end
        end
      endcase
    end
  end

  assign ap_idle = (tapa_state == 2'b00);
  assign ap_done = ap_done__q0;
  assign ap_ready = ap_done__q0;
  assign ap_start__q0 = ap_start;
  assign ap_done__q0 = (tapa_state == 2'b10);

endmodule

